module SCOREBOARD2
(
	input clk,
	input rst,
	input [10:0]row,
	input [10:0]col,
	input [3:0] scoreboard2,
	output reg score_2
);


reg [49:0] s1,s2,s3,s4,s5,s6,s7,s8,s9,s10;
reg [49:0] s11,s12,s13,s14,s15,s16,s17,s18,s19,s20;
reg [49:0] s21,s22,s23,s24,s25,s26,s27,s28,s29,s30;
reg [49:0] s31,s32,s33,s34,s35,s36,s37,s38,s39,s40;
reg [49:0] s41,s42,s43,s44,s45,s46,s47,s48,s49,s50;

wire count;

always@(posedge count)begin
	case(count)
		0:begin
			if(scoreboard2==0)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000111;
				s5 <=50'b11100000000000000000000000000000000000000000000111;
				s6 <=50'b11100000000000000000000000000000000000000000000111;
				s7 <=50'b11100000000000000000000000000000000000000000000111;
				s8 <=50'b11100000000000000000000000000000000000000000000111;
				s9 <=50'b11100000000000000000000000000000000000000000000111;
				s10<=50'b11100000000000000000000000000000000000000000000111;
				s11<=50'b11100000000000000000000000000000000000000000000111;
				s12<=50'b11100000000000000000000000000000000000000000000111;
				s13<=50'b11100000000000000000000000000000000000000000000111;
				s14<=50'b11100000000000000000000000000000000000000000000111;
				s15<=50'b11100000000000000000000000000000000000000000000111;
				s16<=50'b11100000000000000000000000000000000000000000000111;
				s17<=50'b11100000000000000000000000000000000000000000000111;
				s18<=50'b11100000000000000000000000000000000000000000000111;
				s19<=50'b11100000000000000000000000000000000000000000000111;
				s20<=50'b11100000000000000000000000000000000000000000000111;
				s21<=50'b11100000000000000000000000000000000000000000000111;
				s22<=50'b11100000000000000000000000000000000000000000000111;
				s23<=50'b11100000000000000000000000000000000000000000000111;
				s24<=50'b11100000000000000000000000000000000000000000000111;
				s25<=50'b11100000000000000000000000000000000000000000000111;
				s26<=50'b11100000000000000000000000000000000000000000000111;
				s27<=50'b11100000000000000000000000000000000000000000000111;
				s28<=50'b11100000000000000000000000000000000000000000000111;
				s29<=50'b11100000000000000000000000000000000000000000000111;
				s30<=50'b11100000000000000000000000000000000000000000000111;
				s31<=50'b11100000000000000000000000000000000000000000000111;
				s32<=50'b11100000000000000000000000000000000000000000000111;
				s33<=50'b11100000000000000000000000000000000000000000000111;
				s34<=50'b11100000000000000000000000000000000000000000000111;
				s35<=50'b11100000000000000000000000000000000000000000000111;
				s36<=50'b11100000000000000000000000000000000000000000000111;
				s37<=50'b11100000000000000000000000000000000000000000000111;
				s38<=50'b11100000000000000000000000000000000000000000000111;
				s39<=50'b11100000000000000000000000000000000000000000000111;
				s40<=50'b11100000000000000000000000000000000000000000000111;
				s41<=50'b11100000000000000000000000000000000000000000000111;
				s42<=50'b11100000000000000000000000000000000000000000000111;
				s43<=50'b11100000000000000000000000000000000000000000000111;
				s44<=50'b11100000000000000000000000000000000000000000000111;
				s45<=50'b11100000000000000000000000000000000000000000000111;
				s46<=50'b11100000000000000000000000000000000000000000000111;
				s47<=50'b11100000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;				
			end
			
			else if(scoreboard2==1)
			begin
				s1 <=50'b00000000000000000000000000000000000000000000000111;
				s2 <=50'b00000000000000000000000000000000000000000000000111;
				s3 <=50'b00000000000000000000000000000000000000000000000111;
				s4 <=50'b00000000000000000000000000000000000000000000000111;
				s5 <=50'b00000000000000000000000000000000000000000000000111;
				s6 <=50'b00000000000000000000000000000000000000000000000111;
				s7 <=50'b00000000000000000000000000000000000000000000000111;
				s8 <=50'b00000000000000000000000000000000000000000000000111;
				s9 <=50'b00000000000000000000000000000000000000000000000111;
				s10<=50'b00000000000000000000000000000000000000000000000111;
				s11<=50'b00000000000000000000000000000000000000000000000111;
				s12<=50'b00000000000000000000000000000000000000000000000111;
				s13<=50'b00000000000000000000000000000000000000000000000111;
				s14<=50'b00000000000000000000000000000000000000000000000111;
				s15<=50'b00000000000000000000000000000000000000000000000111;
				s16<=50'b00000000000000000000000000000000000000000000000111;
				s17<=50'b00000000000000000000000000000000000000000000000111;
				s18<=50'b00000000000000000000000000000000000000000000000111;
				s19<=50'b00000000000000000000000000000000000000000000000111;
				s20<=50'b00000000000000000000000000000000000000000000000111;
				s21<=50'b00000000000000000000000000000000000000000000000111;
				s22<=50'b00000000000000000000000000000000000000000000000111;
				s23<=50'b00000000000000000000000000000000000000000000000111;
				s24<=50'b00000000000000000000000000000000000000000000000111;
				s25<=50'b00000000000000000000000000000000000000000000000111;
				s26<=50'b00000000000000000000000000000000000000000000000111;
				s27<=50'b00000000000000000000000000000000000000000000000111;
				s28<=50'b00000000000000000000000000000000000000000000000111;
				s29<=50'b00000000000000000000000000000000000000000000000111;
				s30<=50'b00000000000000000000000000000000000000000000000111;
				s31<=50'b00000000000000000000000000000000000000000000000111;
				s32<=50'b00000000000000000000000000000000000000000000000111;
				s33<=50'b00000000000000000000000000000000000000000000000111;
				s34<=50'b00000000000000000000000000000000000000000000000111;
				s35<=50'b00000000000000000000000000000000000000000000000111;
				s36<=50'b00000000000000000000000000000000000000000000000111;
				s37<=50'b00000000000000000000000000000000000000000000000111;
				s38<=50'b00000000000000000000000000000000000000000000000111;
				s39<=50'b00000000000000000000000000000000000000000000000111;
				s40<=50'b00000000000000000000000000000000000000000000000111;
				s41<=50'b00000000000000000000000000000000000000000000000111;
				s42<=50'b00000000000000000000000000000000000000000000000111;
				s43<=50'b00000000000000000000000000000000000000000000000111;
				s44<=50'b00000000000000000000000000000000000000000000000111;
				s45<=50'b00000000000000000000000000000000000000000000000111;
				s46<=50'b00000000000000000000000000000000000000000000000111;
				s47<=50'b00000000000000000000000000000000000000000000000111;
				s48<=50'b00000000000000000000000000000000000000000000000111;
				s49<=50'b00000000000000000000000000000000000000000000000111;
				s50<=50'b00000000000000000000000000000000000000000000000111;				
			end
			
			else if(scoreboard2==2)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b00000000000000000000000000000000000000000000000111;
				s5 <=50'b00000000000000000000000000000000000000000000000111;
				s6 <=50'b00000000000000000000000000000000000000000000000111;
				s7 <=50'b00000000000000000000000000000000000000000000000111;
				s8 <=50'b00000000000000000000000000000000000000000000000111;
				s9 <=50'b00000000000000000000000000000000000000000000000111;
				s10<=50'b00000000000000000000000000000000000000000000000111;
				s11<=50'b00000000000000000000000000000000000000000000000111;
				s12<=50'b00000000000000000000000000000000000000000000000111;
				s13<=50'b00000000000000000000000000000000000000000000000111;
				s14<=50'b00000000000000000000000000000000000000000000000111;
				s15<=50'b00000000000000000000000000000000000000000000000111;
				s16<=50'b00000000000000000000000000000000000000000000000111;
				s17<=50'b00000000000000000000000000000000000000000000000111;
				s18<=50'b00000000000000000000000000000000000000000000000111;
				s19<=50'b00000000000000000000000000000000000000000000000111;
				s20<=50'b00000000000000000000000000000000000000000000000111;
				s21<=50'b00000000000000000000000000000000000000000000000111;
				s22<=50'b00000000000000000000000000000000000000000000000111;
				s23<=50'b00000000000000000000000000000000000000000000000111;
				s24<=50'b00000000000000000000000000000000000000000000000111;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b11100000000000000000000000000000000000000000000000;
				s28<=50'b11100000000000000000000000000000000000000000000000;
				s29<=50'b11100000000000000000000000000000000000000000000000;
				s30<=50'b11100000000000000000000000000000000000000000000000;
				s31<=50'b11100000000000000000000000000000000000000000000000;
				s32<=50'b11100000000000000000000000000000000000000000000000;
				s33<=50'b11100000000000000000000000000000000000000000000000;
				s34<=50'b11100000000000000000000000000000000000000000000000;
				s35<=50'b11100000000000000000000000000000000000000000000000;
				s36<=50'b11100000000000000000000000000000000000000000000000;
				s37<=50'b11100000000000000000000000000000000000000000000000;
				s38<=50'b11100000000000000000000000000000000000000000000000;
				s39<=50'b11100000000000000000000000000000000000000000000000;
				s40<=50'b11100000000000000000000000000000000000000000000000;
				s41<=50'b11100000000000000000000000000000000000000000000000;
				s42<=50'b11100000000000000000000000000000000000000000000000;
				s43<=50'b11100000000000000000000000000000000000000000000000;
				s44<=50'b11100000000000000000000000000000000000000000000000;
				s45<=50'b11100000000000000000000000000000000000000000000000;
				s46<=50'b11100000000000000000000000000000000000000000000000;
				s47<=50'b11100000000000000000000000000000000000000000000000;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;				
			end
			
			else if(scoreboard2==3)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b00000000000000000000000000000000000000000000000111;
				s5 <=50'b00000000000000000000000000000000000000000000000111;
				s6 <=50'b00000000000000000000000000000000000000000000000111;
				s7 <=50'b00000000000000000000000000000000000000000000000111;
				s8 <=50'b00000000000000000000000000000000000000000000000111;
				s9 <=50'b00000000000000000000000000000000000000000000000111;
				s10<=50'b00000000000000000000000000000000000000000000000111;
				s11<=50'b00000000000000000000000000000000000000000000000111;
				s12<=50'b00000000000000000000000000000000000000000000000111;
				s13<=50'b00000000000000000000000000000000000000000000000111;
				s14<=50'b00000000000000000000000000000000000000000000000111;
				s15<=50'b00000000000000000000000000000000000000000000000111;
				s16<=50'b00000000000000000000000000000000000000000000000111;
				s17<=50'b00000000000000000000000000000000000000000000000111;
				s18<=50'b00000000000000000000000000000000000000000000000111;
				s19<=50'b00000000000000000000000000000000000000000000000111;
				s20<=50'b00000000000000000000000000000000000000000000000111;
				s21<=50'b00000000000000000000000000000000000000000000000111;
				s22<=50'b00000000000000000000000000000000000000000000000111;
				s23<=50'b00000000000000000000000000000000000000000000000111;
				s24<=50'b00000000000000000000000000000000000000000000000111;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b00000000000000000000000000000000000000000000000111;
				s28<=50'b00000000000000000000000000000000000000000000000111;
				s29<=50'b00000000000000000000000000000000000000000000000111;
				s30<=50'b00000000000000000000000000000000000000000000000111;
				s31<=50'b00000000000000000000000000000000000000000000000111;
				s32<=50'b00000000000000000000000000000000000000000000000111;
				s33<=50'b00000000000000000000000000000000000000000000000111;
				s34<=50'b00000000000000000000000000000000000000000000000111;
				s35<=50'b00000000000000000000000000000000000000000000000111;
				s36<=50'b00000000000000000000000000000000000000000000000111;
				s37<=50'b00000000000000000000000000000000000000000000000111;
				s38<=50'b00000000000000000000000000000000000000000000000111;
				s39<=50'b00000000000000000000000000000000000000000000000111;
				s40<=50'b00000000000000000000000000000000000000000000000111;
				s41<=50'b00000000000000000000000000000000000000000000000111;
				s42<=50'b00000000000000000000000000000000000000000000000111;
				s43<=50'b00000000000000000000000000000000000000000000000111;
				s44<=50'b00000000000000000000000000000000000000000000000111;
				s45<=50'b00000000000000000000000000000000000000000000000111;
				s46<=50'b00000000000000000000000000000000000000000000000111;
				s47<=50'b00000000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;				
			end
			
			else if(scoreboard2==4)
			begin
				s1 <=50'b11100000000000000000000000000000000000000000000000;
				s2 <=50'b11100000000000000000000000000000000000000000000000;
				s3 <=50'b11100000000000000000000000000000000000000000000000;
				s4 <=50'b11100000000000000000000000000000000000000000000000;
				s5 <=50'b11100000000000000000000000000000000000000000000000;
				s6 <=50'b11100000000000000000000000000000000000000000000000;
				s7 <=50'b11100000000000000000000000000000000000000000000000;
				s8 <=50'b11100000000000000000000000000000000000000000000000;
				s9 <=50'b11100000000000000000000000000000000000000000000000;
				s10<=50'b11100000000000000000000000000000000000000000000000;
				s11<=50'b11100000000000000000000000000000000000000000000000;
				s12<=50'b11100000000000000000000000000000000000000000000000;
				s13<=50'b11100000000000000000000000000000000000000000000000;
				s14<=50'b11100000000000000000000000000000000000000000000000;
				s15<=50'b11100000000000000000000000000000000000000000000000;
				s16<=50'b11100000000000000000001110000000000000000000000000;
				s17<=50'b11100000000000000000001110000000000000000000000000;
				s18<=50'b11100000000000000000001110000000000000000000000000;
				s19<=50'b11100000000000000000001110000000000000000000000000;
				s20<=50'b11100000000000000000001110000000000000000000000000;
				s21<=50'b11100000000000000000001110000000000000000000000000;
				s22<=50'b11100000000000000000001110000000000000000000000000;
				s23<=50'b11100000000000000000001110000000000000000000000000;
				s24<=50'b11100000000000000000001110000000000000000000000000;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b00000000000000000000001110000000000000000000000000;
				s28<=50'b00000000000000000000001110000000000000000000000000;
				s29<=50'b00000000000000000000001110000000000000000000000000;
				s30<=50'b00000000000000000000001110000000000000000000000000;
				s31<=50'b00000000000000000000001110000000000000000000000000;
				s32<=50'b00000000000000000000001110000000000000000000000000;
				s33<=50'b00000000000000000000001110000000000000000000000000;
				s34<=50'b00000000000000000000001110000000000000000000000000;
				s35<=50'b00000000000000000000001110000000000000000000000000;
				s36<=50'b00000000000000000000001110000000000000000000000000;
				s37<=50'b00000000000000000000001110000000000000000000000000;
				s38<=50'b00000000000000000000001110000000000000000000000000;
				s39<=50'b00000000000000000000001110000000000000000000000000;
				s40<=50'b00000000000000000000001110000000000000000000000000;
				s41<=50'b00000000000000000000001110000000000000000000000000;
				s42<=50'b00000000000000000000001110000000000000000000000000;
				s43<=50'b00000000000000000000001110000000000000000000000000;
				s44<=50'b00000000000000000000001110000000000000000000000000;
				s45<=50'b00000000000000000000001110000000000000000000000000;
				s46<=50'b00000000000000000000001110000000000000000000000000;
				s47<=50'b00000000000000000000001110000000000000000000000000;
				s48<=50'b00000000000000000000001110000000000000000000000000;
				s49<=50'b00000000000000000000001110000000000000000000000000;
				s50<=50'b00000000000000000000001110000000000000000000000000;				
			end
			
			else if(scoreboard2==5)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000000;
				s5 <=50'b11100000000000000000000000000000000000000000000000;
				s6 <=50'b11100000000000000000000000000000000000000000000000;
				s7 <=50'b11100000000000000000000000000000000000000000000000;
				s8 <=50'b11100000000000000000000000000000000000000000000000;
				s9 <=50'b11100000000000000000000000000000000000000000000000;
				s10<=50'b11100000000000000000000000000000000000000000000000;
				s11<=50'b11100000000000000000000000000000000000000000000000;
				s12<=50'b11100000000000000000000000000000000000000000000000;
				s13<=50'b11100000000000000000000000000000000000000000000000;
				s14<=50'b11100000000000000000000000000000000000000000000000;
				s15<=50'b11100000000000000000000000000000000000000000000000;
				s16<=50'b11100000000000000000000000000000000000000000000000;
				s17<=50'b11100000000000000000000000000000000000000000000000;
				s18<=50'b11100000000000000000000000000000000000000000000000;
				s19<=50'b11100000000000000000000000000000000000000000000000;
				s20<=50'b11100000000000000000000000000000000000000000000000;
				s21<=50'b11100000000000000000000000000000000000000000000000;
				s22<=50'b11100000000000000000000000000000000000000000000000;
				s23<=50'b11100000000000000000000000000000000000000000000000;
				s24<=50'b11100000000000000000000000000000000000000000000000;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b00000000000000000000000000000000000000000000000111;
				s28<=50'b00000000000000000000000000000000000000000000000111;
				s29<=50'b00000000000000000000000000000000000000000000000111;
				s30<=50'b00000000000000000000000000000000000000000000000111;
				s31<=50'b00000000000000000000000000000000000000000000000111;
				s32<=50'b00000000000000000000000000000000000000000000000111;
				s33<=50'b00000000000000000000000000000000000000000000000111;
				s34<=50'b00000000000000000000000000000000000000000000000111;
				s35<=50'b00000000000000000000000000000000000000000000000111;
				s36<=50'b00000000000000000000000000000000000000000000000111;
				s37<=50'b00000000000000000000000000000000000000000000000111;
				s38<=50'b00000000000000000000000000000000000000000000000111;
				s39<=50'b00000000000000000000000000000000000000000000000111;
				s40<=50'b00000000000000000000000000000000000000000000000111;
				s41<=50'b00000000000000000000000000000000000000000000000111;
				s42<=50'b00000000000000000000000000000000000000000000000111;
				s43<=50'b00000000000000000000000000000000000000000000000111;
				s44<=50'b00000000000000000000000000000000000000000000000111;
				s45<=50'b00000000000000000000000000000000000000000000000111;
				s46<=50'b00000000000000000000000000000000000000000000000111;
				s47<=50'b00000000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;			
			end
			
			else if(scoreboard2==6)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000000;
				s5 <=50'b11100000000000000000000000000000000000000000000000;
				s6 <=50'b11100000000000000000000000000000000000000000000000;
				s7 <=50'b11100000000000000000000000000000000000000000000000;
				s8 <=50'b11100000000000000000000000000000000000000000000000;
				s9 <=50'b11100000000000000000000000000000000000000000000000;
				s10<=50'b11100000000000000000000000000000000000000000000000;
				s11<=50'b11100000000000000000000000000000000000000000000000;
				s12<=50'b11100000000000000000000000000000000000000000000000;
				s13<=50'b11100000000000000000000000000000000000000000000000;
				s14<=50'b11100000000000000000000000000000000000000000000000;
				s15<=50'b11100000000000000000000000000000000000000000000000;
				s16<=50'b11100000000000000000000000000000000000000000000000;
				s17<=50'b11100000000000000000000000000000000000000000000000;
				s18<=50'b11100000000000000000000000000000000000000000000000;
				s19<=50'b11100000000000000000000000000000000000000000000000;
				s20<=50'b11100000000000000000000000000000000000000000000000;
				s21<=50'b11100000000000000000000000000000000000000000000000;
				s22<=50'b11100000000000000000000000000000000000000000000000;
				s23<=50'b11100000000000000000000000000000000000000000000000;
				s24<=50'b11100000000000000000000000000000000000000000000000;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b11100000000000000000000000000000000000000000000111;
				s28<=50'b11100000000000000000000000000000000000000000000111;
				s29<=50'b11100000000000000000000000000000000000000000000111;
				s30<=50'b11100000000000000000000000000000000000000000000111;
				s31<=50'b11100000000000000000000000000000000000000000000111;
				s32<=50'b11100000000000000000000000000000000000000000000111;
				s33<=50'b11100000000000000000000000000000000000000000000111;
				s34<=50'b11100000000000000000000000000000000000000000000111;
				s35<=50'b11100000000000000000000000000000000000000000000111;
				s36<=50'b11100000000000000000000000000000000000000000000111;
				s37<=50'b11100000000000000000000000000000000000000000000111;
				s38<=50'b11100000000000000000000000000000000000000000000111;
				s39<=50'b11100000000000000000000000000000000000000000000111;
				s40<=50'b11100000000000000000000000000000000000000000000111;
				s41<=50'b11100000000000000000000000000000000000000000000111;
				s42<=50'b11100000000000000000000000000000000000000000000111;
				s43<=50'b11100000000000000000000000000000000000000000000111;
				s44<=50'b11100000000000000000000000000000000000000000000111;
				s45<=50'b11100000000000000000000000000000000000000000000111;
				s46<=50'b11100000000000000000000000000000000000000000000111;
				s47<=50'b11100000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;
			end
			
			else if(scoreboard2==7)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b00000000000000000000000000000000000000000000000111;
				s5 <=50'b00000000000000000000000000000000000000000000000111;
				s6 <=50'b00000000000000000000000000000000000000000000000111;
				s7 <=50'b00000000000000000000000000000000000000000000000111;
				s8 <=50'b00000000000000000000000000000000000000000000000111;
				s9 <=50'b00000000000000000000000000000000000000000000000111;
				s10<=50'b00000000000000000000000000000000000000000000000111;
				s11<=50'b00000000000000000000000000000000000000000000000111;
				s12<=50'b00000000000000000000000000000000000000000000000111;
				s13<=50'b00000000000000000000000000000000000000000000000111;
				s14<=50'b00000000000000000000000000000000000000000000000111;
				s15<=50'b00000000000000000000000000000000000000000000000111;
				s16<=50'b00000000000000000000000000000000000000000000000111;
				s17<=50'b00000000000000000000000000000000000000000000000111;
				s18<=50'b00000000000000000000000000000000000000000000000111;
				s19<=50'b00000000000000000000000000000000000000000000000111;
				s20<=50'b00000000000000000000000000000000000000000000000111;
				s21<=50'b00000000000000000000000000000000000000000000000111;
				s22<=50'b00000000000000000000000000000000000000000000000111;
				s23<=50'b00000000000000000000000000000000000000000000000111;
				s24<=50'b00000000000000000000000000000000000000000000000111;
				s25<=50'b00000000000000000000000000000000000000000000000111;
				s26<=50'b00000000000000000000000000000000000000000000000111;
				s27<=50'b00000000000000000000000000000000000000000000000111;
				s28<=50'b00000000000000000000000000000000000000000000000111;
				s29<=50'b00000000000000000000000000000000000000000000000111;
				s30<=50'b00000000000000000000000000000000000000000000000111;
				s31<=50'b00000000000000000000000000000000000000000000000111;
				s32<=50'b00000000000000000000000000000000000000000000000111;
				s33<=50'b00000000000000000000000000000000000000000000000111;
				s34<=50'b00000000000000000000000000000000000000000000000111;
				s35<=50'b00000000000000000000000000000000000000000000000111;
				s36<=50'b00000000000000000000000000000000000000000000000111;
				s37<=50'b00000000000000000000000000000000000000000000000111;
				s38<=50'b00000000000000000000000000000000000000000000000111;
				s39<=50'b00000000000000000000000000000000000000000000000111;
				s40<=50'b00000000000000000000000000000000000000000000000111;
				s41<=50'b00000000000000000000000000000000000000000000000111;
				s42<=50'b00000000000000000000000000000000000000000000000111;
				s43<=50'b00000000000000000000000000000000000000000000000111;
				s44<=50'b00000000000000000000000000000000000000000000000111;
				s45<=50'b00000000000000000000000000000000000000000000000111;
				s46<=50'b00000000000000000000000000000000000000000000000111;
				s47<=50'b00000000000000000000000000000000000000000000000111;
				s48<=50'b00000000000000000000000000000000000000000000000111;
				s49<=50'b00000000000000000000000000000000000000000000000111;
				s50<=50'b00000000000000000000000000000000000000000000000111;				
			end
			
			else if(scoreboard2==8)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000111;
				s5 <=50'b11100000000000000000000000000000000000000000000111;
				s6 <=50'b11100000000000000000000000000000000000000000000111;
				s7 <=50'b11100000000000000000000000000000000000000000000111;
				s8 <=50'b11100000000000000000000000000000000000000000000111;
				s9 <=50'b11100000000000000000000000000000000000000000000111;
				s10<=50'b11100000000000000000000000000000000000000000000111;
				s11<=50'b11100000000000000000000000000000000000000000000111;
				s12<=50'b11100000000000000000000000000000000000000000000111;
				s13<=50'b11100000000000000000000000000000000000000000000111;
				s14<=50'b11100000000000000000000000000000000000000000000111;
				s15<=50'b11100000000000000000000000000000000000000000000111;
				s16<=50'b11100000000000000000000000000000000000000000000111;
				s17<=50'b11100000000000000000000000000000000000000000000111;
				s18<=50'b11100000000000000000000000000000000000000000000111;
				s19<=50'b11100000000000000000000000000000000000000000000111;
				s20<=50'b11100000000000000000000000000000000000000000000111;
				s21<=50'b11100000000000000000000000000000000000000000000111;
				s22<=50'b11100000000000000000000000000000000000000000000111;
				s23<=50'b11100000000000000000000000000000000000000000000111;
				s24<=50'b11100000000000000000000000000000000000000000000111;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b11100000000000000000000000000000000000000000000111;
				s28<=50'b11100000000000000000000000000000000000000000000111;
				s29<=50'b11100000000000000000000000000000000000000000000111;
				s30<=50'b11100000000000000000000000000000000000000000000111;
				s31<=50'b11100000000000000000000000000000000000000000000111;
				s32<=50'b11100000000000000000000000000000000000000000000111;
				s33<=50'b11100000000000000000000000000000000000000000000111;
				s34<=50'b11100000000000000000000000000000000000000000000111;
				s35<=50'b11100000000000000000000000000000000000000000000111;
				s36<=50'b11100000000000000000000000000000000000000000000111;
				s37<=50'b11100000000000000000000000000000000000000000000111;
				s38<=50'b11100000000000000000000000000000000000000000000111;
				s39<=50'b11100000000000000000000000000000000000000000000111;
				s40<=50'b11100000000000000000000000000000000000000000000111;
				s41<=50'b11100000000000000000000000000000000000000000000111;
				s42<=50'b11100000000000000000000000000000000000000000000111;
				s43<=50'b11100000000000000000000000000000000000000000000111;
				s44<=50'b11100000000000000000000000000000000000000000000111;
				s45<=50'b11100000000000000000000000000000000000000000000111;
				s46<=50'b11100000000000000000000000000000000000000000000111;
				s47<=50'b11100000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;					
			end
			
			else if(scoreboard2==9)
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000111;
				s5 <=50'b11100000000000000000000000000000000000000000000111;
				s6 <=50'b11100000000000000000000000000000000000000000000111;
				s7 <=50'b11100000000000000000000000000000000000000000000111;
				s8 <=50'b11100000000000000000000000000000000000000000000111;
				s9 <=50'b11100000000000000000000000000000000000000000000111;
				s10<=50'b11100000000000000000000000000000000000000000000111;
				s11<=50'b11100000000000000000000000000000000000000000000111;
				s12<=50'b11100000000000000000000000000000000000000000000111;
				s13<=50'b11100000000000000000000000000000000000000000000111;
				s14<=50'b11100000000000000000000000000000000000000000000111;
				s15<=50'b11100000000000000000000000000000000000000000000111;
				s16<=50'b11100000000000000000000000000000000000000000000111;
				s17<=50'b11100000000000000000000000000000000000000000000111;
				s18<=50'b11100000000000000000000000000000000000000000000111;
				s19<=50'b11100000000000000000000000000000000000000000000111;
				s20<=50'b11100000000000000000000000000000000000000000000111;
				s21<=50'b11100000000000000000000000000000000000000000000111;
				s22<=50'b11100000000000000000000000000000000000000000000111;
				s23<=50'b11100000000000000000000000000000000000000000000111;
				s24<=50'b11100000000000000000000000000000000000000000000111;
				s25<=50'b11111111111111111111111111111111111111111111111111;
				s26<=50'b11111111111111111111111111111111111111111111111111;
				s27<=50'b00000000000000000000000000000000000000000000000111;
				s28<=50'b00000000000000000000000000000000000000000000000111;
				s29<=50'b00000000000000000000000000000000000000000000000111;
				s30<=50'b00000000000000000000000000000000000000000000000111;
				s31<=50'b00000000000000000000000000000000000000000000000111;
				s32<=50'b00000000000000000000000000000000000000000000000111;
				s33<=50'b00000000000000000000000000000000000000000000000111;
				s34<=50'b00000000000000000000000000000000000000000000000111;
				s35<=50'b00000000000000000000000000000000000000000000000111;
				s36<=50'b00000000000000000000000000000000000000000000000111;
				s37<=50'b00000000000000000000000000000000000000000000000111;
				s38<=50'b00000000000000000000000000000000000000000000000111;
				s39<=50'b00000000000000000000000000000000000000000000000111;
				s40<=50'b00000000000000000000000000000000000000000000000111;
				s41<=50'b00000000000000000000000000000000000000000000000111;
				s42<=50'b00000000000000000000000000000000000000000000000111;
				s43<=50'b00000000000000000000000000000000000000000000000111;
				s44<=50'b00000000000000000000000000000000000000000000000111;
				s45<=50'b00000000000000000000000000000000000000000000000111;
				s46<=50'b00000000000000000000000000000000000000000000000111;
				s47<=50'b00000000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;				
			end	
		
		else
			begin
				s1 <=50'b11111111111111111111111111111111111111111111111111;
				s2 <=50'b11111111111111111111111111111111111111111111111111;
				s3 <=50'b11111111111111111111111111111111111111111111111111;
				s4 <=50'b11100000000000000000000000000000000000000000000111;
				s5 <=50'b11100000000000000000000000000000000000000000000111;
				s6 <=50'b11100000000000000000000000000000000000000000000111;
				s7 <=50'b11100000000000000000000000000000000000000000000111;
				s8 <=50'b11100000000000000000000000000000000000000000000111;
				s9 <=50'b11100000000000000000000000000000000000000000000111;
				s10<=50'b11100000000000000000000000000000000000000000000111;
				s11<=50'b11100000000000000000000000000000000000000000000111;
				s12<=50'b11100000000000000000000000000000000000000000000111;
				s13<=50'b11100000000000000000000000000000000000000000000111;
				s14<=50'b11100000000000000000000000000000000000000000000111;
				s15<=50'b11100000000000000000000000000000000000000000000111;
				s16<=50'b11100000000000000000000000000000000000000000000111;
				s17<=50'b11100000000000000000000000000000000000000000000111;
				s18<=50'b11100000000000000000000000000000000000000000000111;
				s19<=50'b11100000000000000000000000000000000000000000000111;
				s20<=50'b11100000000000000000000000000000000000000000000111;
				s21<=50'b11100000000000000000000000000000000000000000000111;
				s22<=50'b11100000000000000000000000000000000000000000000111;
				s23<=50'b11100000000000000000000000000000000000000000000111;
				s24<=50'b11100000000000000000000000000000000000000000000111;
				s25<=50'b11100000000000000000000000000000000000000000000111;
				s26<=50'b11100000000000000000000000000000000000000000000111;
				s27<=50'b11100000000000000000000000000000000000000000000111;
				s28<=50'b11100000000000000000000000000000000000000000000111;
				s29<=50'b11100000000000000000000000000000000000000000000111;
				s30<=50'b11100000000000000000000000000000000000000000000111;
				s31<=50'b11100000000000000000000000000000000000000000000111;
				s32<=50'b11100000000000000000000000000000000000000000000111;
				s33<=50'b11100000000000000000000000000000000000000000000111;
				s34<=50'b11100000000000000000000000000000000000000000000111;
				s35<=50'b11100000000000000000000000000000000000000000000111;
				s36<=50'b11100000000000000000000000000000000000000000000111;
				s37<=50'b11100000000000000000000000000000000000000000000111;
				s38<=50'b11100000000000000000000000000000000000000000000111;
				s39<=50'b11100000000000000000000000000000000000000000000111;
				s40<=50'b11100000000000000000000000000000000000000000000111;
				s41<=50'b11100000000000000000000000000000000000000000000111;
				s42<=50'b11100000000000000000000000000000000000000000000111;
				s43<=50'b11100000000000000000000000000000000000000000000111;
				s44<=50'b11100000000000000000000000000000000000000000000111;
				s45<=50'b11100000000000000000000000000000000000000000000111;
				s46<=50'b11100000000000000000000000000000000000000000000111;
				s47<=50'b11100000000000000000000000000000000000000000000111;
				s48<=50'b11111111111111111111111111111111111111111111111111;
				s49<=50'b11111111111111111111111111111111111111111111111111;
				s50<=50'b11111111111111111111111111111111111111111111111111;				
			end
		end
	endcase		
end

always@(posedge clk)begin
	case(row)
				600: begin
						case(col)
							730:score_2<=s50[49];
							731:score_2<=s50[48];
							732:score_2<=s50[47];
							733:score_2<=s50[46];
							734:score_2<=s50[45];
							735:score_2<=s50[44];
							736:score_2<=s50[43];
							737:score_2<=s50[42];
							738:score_2<=s50[41];
							739:score_2<=s50[40];
							740:score_2<=s50[39];
							741:score_2<=s50[38];
							742:score_2<=s50[37];
							743:score_2<=s50[36];
							744:score_2<=s50[35];
							745:score_2<=s50[34];
							746:score_2<=s50[33];
							747:score_2<=s50[32];
							748:score_2<=s50[31];
							749:score_2<=s50[30];
							750:score_2<=s50[29];
							751:score_2<=s50[28];
							752:score_2<=s50[27];
							753:score_2<=s50[26];
							754:score_2<=s50[25];
							755:score_2<=s50[24];
							756:score_2<=s50[23];
							757:score_2<=s50[22];
							758:score_2<=s50[21];
							759:score_2<=s50[20];
							760:score_2<=s50[19];
							761:score_2<=s50[18];
							762:score_2<=s50[17];
							763:score_2<=s50[16];
							764:score_2<=s50[15];
							765:score_2<=s50[14];
							766:score_2<=s50[13];
							767:score_2<=s50[12];
							768:score_2<=s50[11];
							769:score_2<=s50[10];
							770:score_2<=s50[9];
							771:score_2<=s50[8];
							772:score_2<=s50[7];
							773:score_2<=s50[6];
							774:score_2<=s50[5];
							775:score_2<=s50[4];
							776:score_2<=s50[3];
							777:score_2<=s50[2];
							778:score_2<=s50[1];
							779:score_2<=s50[0];
							default:score_2<=0;
						endcase
					end
					599: begin
						case(col)
							730:score_2<=s49[49];
							731:score_2<=s49[48];
							732:score_2<=s49[47];
							733:score_2<=s49[46];
							734:score_2<=s49[45];
							735:score_2<=s49[44];
							736:score_2<=s49[43];
							737:score_2<=s49[42];
							738:score_2<=s49[41];
							739:score_2<=s49[40];
							740:score_2<=s49[39];
							741:score_2<=s49[38];
							742:score_2<=s49[37];
							743:score_2<=s49[36];
							744:score_2<=s49[35];
							745:score_2<=s49[34];
							746:score_2<=s49[33];
							747:score_2<=s49[32];
							748:score_2<=s49[31];
							749:score_2<=s49[30];
							750:score_2<=s49[29];
							751:score_2<=s49[28];
							752:score_2<=s49[27];
							753:score_2<=s49[26];
							754:score_2<=s49[25];
							755:score_2<=s49[24];
							756:score_2<=s49[23];
							757:score_2<=s49[22];
							758:score_2<=s49[21];
							759:score_2<=s49[20];
							760:score_2<=s49[19];
							761:score_2<=s49[18];
							762:score_2<=s49[17];
							763:score_2<=s49[16];
							764:score_2<=s49[15];
							765:score_2<=s49[14];
							766:score_2<=s49[13];
							767:score_2<=s49[12];
							768:score_2<=s49[11];
							769:score_2<=s49[10];
							770:score_2<=s49[9];
							771:score_2<=s49[8];
							772:score_2<=s49[7];
							773:score_2<=s49[6];
							774:score_2<=s49[5];
							775:score_2<=s49[4];
							776:score_2<=s49[3];
							777:score_2<=s49[2];
							778:score_2<=s49[1];
							779:score_2<=s49[0];
							default:score_2<=0;
						endcase
					end
					598: begin
						case(col)
							730:score_2<=s48[49];
							731:score_2<=s48[48];
							732:score_2<=s48[47];
							733:score_2<=s48[46];
							734:score_2<=s48[45];
							735:score_2<=s48[44];
							736:score_2<=s48[43];
							737:score_2<=s48[42];
							738:score_2<=s48[41];
							739:score_2<=s48[40];
							740:score_2<=s48[39];
							741:score_2<=s48[38];
							742:score_2<=s48[37];
							743:score_2<=s48[36];
							744:score_2<=s48[35];
							745:score_2<=s48[34];
							746:score_2<=s48[33];
							747:score_2<=s48[32];
							748:score_2<=s48[31];
							749:score_2<=s48[30];
							750:score_2<=s48[29];
							751:score_2<=s48[28];
							752:score_2<=s48[27];
							753:score_2<=s48[26];
							754:score_2<=s48[25];
							755:score_2<=s48[24];
							756:score_2<=s48[23];
							757:score_2<=s48[22];
							758:score_2<=s48[21];
							759:score_2<=s48[20];
							760:score_2<=s48[19];
							761:score_2<=s48[18];
							762:score_2<=s48[17];
							763:score_2<=s48[16];
							764:score_2<=s48[15];
							765:score_2<=s48[14];
							766:score_2<=s48[13];
							767:score_2<=s48[12];
							768:score_2<=s48[11];
							769:score_2<=s48[10];
							770:score_2<=s48[9];
							771:score_2<=s48[8];
							772:score_2<=s48[7];
							773:score_2<=s48[6];
							774:score_2<=s48[5];
							775:score_2<=s48[4];
							776:score_2<=s48[3];
							777:score_2<=s48[2];
							778:score_2<=s48[1];
							779:score_2<=s48[0];
							default:score_2<=0;
						endcase
					end
					597: begin
						case(col)
							730:score_2<=s47[49];
							731:score_2<=s47[48];
							732:score_2<=s47[47];
							733:score_2<=s47[46];
							734:score_2<=s47[45];
							735:score_2<=s47[44];
							736:score_2<=s47[43];
							737:score_2<=s47[42];
							738:score_2<=s47[41];
							739:score_2<=s47[40];
							740:score_2<=s47[39];
							741:score_2<=s47[38];
							742:score_2<=s47[37];
							743:score_2<=s47[36];
							744:score_2<=s47[35];
							745:score_2<=s47[34];
							746:score_2<=s47[33];
							747:score_2<=s47[32];
							748:score_2<=s47[31];
							749:score_2<=s47[30];
							750:score_2<=s47[29];
							751:score_2<=s47[28];
							752:score_2<=s47[27];
							753:score_2<=s47[26];
							754:score_2<=s47[25];
							755:score_2<=s47[24];
							756:score_2<=s47[23];
							757:score_2<=s47[22];
							758:score_2<=s47[21];
							759:score_2<=s47[20];
							760:score_2<=s47[19];
							761:score_2<=s47[18];
							762:score_2<=s47[17];
							763:score_2<=s47[16];
							764:score_2<=s47[15];
							765:score_2<=s47[14];
							766:score_2<=s47[13];
							767:score_2<=s47[12];
							768:score_2<=s47[11];
							769:score_2<=s47[10];
							770:score_2<=s47[9];
							771:score_2<=s47[8];
							772:score_2<=s47[7];
							773:score_2<=s47[6];
							774:score_2<=s47[5];
							775:score_2<=s47[4];
							776:score_2<=s47[3];
							777:score_2<=s47[2];
							778:score_2<=s47[1];
							779:score_2<=s47[0];
							default:score_2<=0;
						endcase
					end
					596: begin
						case(col)
							730:score_2<=s46[49];
							731:score_2<=s46[48];
							732:score_2<=s46[47];
							733:score_2<=s46[46];
							734:score_2<=s46[45];
							735:score_2<=s46[44];
							736:score_2<=s46[43];
							737:score_2<=s46[42];
							738:score_2<=s46[41];
							739:score_2<=s46[40];
							740:score_2<=s46[39];
							741:score_2<=s46[38];
							742:score_2<=s46[37];
							743:score_2<=s46[36];
							744:score_2<=s46[35];
							745:score_2<=s46[34];
							746:score_2<=s46[33];
							747:score_2<=s46[32];
							748:score_2<=s46[31];
							749:score_2<=s46[30];
							750:score_2<=s46[29];
							751:score_2<=s46[28];
							752:score_2<=s46[27];
							753:score_2<=s46[26];
							754:score_2<=s46[25];
							755:score_2<=s46[24];
							756:score_2<=s46[23];
							757:score_2<=s46[22];
							758:score_2<=s46[21];
							759:score_2<=s46[20];
							760:score_2<=s46[19];
							761:score_2<=s46[18];
							762:score_2<=s46[17];
							763:score_2<=s46[16];
							764:score_2<=s46[15];
							765:score_2<=s46[14];
							766:score_2<=s46[13];
							767:score_2<=s46[12];
							768:score_2<=s46[11];
							769:score_2<=s46[10];
							770:score_2<=s46[9];
							771:score_2<=s46[8];
							772:score_2<=s46[7];
							773:score_2<=s46[6];
							774:score_2<=s46[5];
							775:score_2<=s46[4];
							776:score_2<=s46[3];
							777:score_2<=s46[2];
							778:score_2<=s46[1];
							779:score_2<=s46[0];
							default:score_2<=0;
						endcase
					end
					595: begin
						case(col)
							730:score_2<=s45[49];
							731:score_2<=s45[48];
							732:score_2<=s45[47];
							733:score_2<=s45[46];
							734:score_2<=s45[45];
							735:score_2<=s45[44];
							736:score_2<=s45[43];
							737:score_2<=s45[42];
							738:score_2<=s45[41];
							739:score_2<=s45[40];
							740:score_2<=s45[39];
							741:score_2<=s45[38];
							742:score_2<=s45[37];
							743:score_2<=s45[36];
							744:score_2<=s45[35];
							745:score_2<=s45[34];
							746:score_2<=s45[33];
							747:score_2<=s45[32];
							748:score_2<=s45[31];
							749:score_2<=s45[30];
							750:score_2<=s45[29];
							751:score_2<=s45[28];
							752:score_2<=s45[27];
							753:score_2<=s45[26];
							754:score_2<=s45[25];
							755:score_2<=s45[24];
							756:score_2<=s45[23];
							757:score_2<=s45[22];
							758:score_2<=s45[21];
							759:score_2<=s45[20];
							760:score_2<=s45[19];
							761:score_2<=s45[18];
							762:score_2<=s45[17];
							763:score_2<=s45[16];
							764:score_2<=s45[15];
							765:score_2<=s45[14];
							766:score_2<=s45[13];
							767:score_2<=s45[12];
							768:score_2<=s45[11];
							769:score_2<=s45[10];
							770:score_2<=s45[9];
							771:score_2<=s45[8];
							772:score_2<=s45[7];
							773:score_2<=s45[6];
							774:score_2<=s45[5];
							775:score_2<=s45[4];
							776:score_2<=s45[3];
							777:score_2<=s45[2];
							778:score_2<=s45[1];
							779:score_2<=s45[0];
							default:score_2<=0;
						endcase
					end
					594: begin
						case(col)
							730:score_2<=s44[49];
							731:score_2<=s44[48];
							732:score_2<=s44[47];
							733:score_2<=s44[46];
							734:score_2<=s44[45];
							735:score_2<=s44[44];
							736:score_2<=s44[43];
							737:score_2<=s44[42];
							738:score_2<=s44[41];
							739:score_2<=s44[40];
							740:score_2<=s44[39];
							741:score_2<=s44[38];
							742:score_2<=s44[37];
							743:score_2<=s44[36];
							744:score_2<=s44[35];
							745:score_2<=s44[34];
							746:score_2<=s44[33];
							747:score_2<=s44[32];
							748:score_2<=s44[31];
							749:score_2<=s44[30];
							750:score_2<=s44[29];
							751:score_2<=s44[28];
							752:score_2<=s44[27];
							753:score_2<=s44[26];
							754:score_2<=s44[25];
							755:score_2<=s44[24];
							756:score_2<=s44[23];
							757:score_2<=s44[22];
							758:score_2<=s44[21];
							759:score_2<=s44[20];
							760:score_2<=s44[19];
							761:score_2<=s44[18];
							762:score_2<=s44[17];
							763:score_2<=s44[16];
							764:score_2<=s44[15];
							765:score_2<=s44[14];
							766:score_2<=s44[13];
							767:score_2<=s44[12];
							768:score_2<=s44[11];
							769:score_2<=s44[10];
							770:score_2<=s44[9];
							771:score_2<=s44[8];
							772:score_2<=s44[7];
							773:score_2<=s44[6];
							774:score_2<=s44[5];
							775:score_2<=s44[4];
							776:score_2<=s44[3];
							777:score_2<=s44[2];
							778:score_2<=s44[1];
							779:score_2<=s44[0];
							default:score_2<=0;
						endcase
					end
					593: begin
						case(col)
							730:score_2<=s43[49];
							731:score_2<=s43[48];
							732:score_2<=s43[47];
							733:score_2<=s43[46];
							734:score_2<=s43[45];
							735:score_2<=s43[44];
							736:score_2<=s43[43];
							737:score_2<=s43[42];
							738:score_2<=s43[41];
							739:score_2<=s43[40];
							740:score_2<=s43[39];
							741:score_2<=s43[38];
							742:score_2<=s43[37];
							743:score_2<=s43[36];
							744:score_2<=s43[35];
							745:score_2<=s43[34];
							746:score_2<=s43[33];
							747:score_2<=s43[32];
							748:score_2<=s43[31];
							749:score_2<=s43[30];
							750:score_2<=s43[29];
							751:score_2<=s43[28];
							752:score_2<=s43[27];
							753:score_2<=s43[26];
							754:score_2<=s43[25];
							755:score_2<=s43[24];
							756:score_2<=s43[23];
							757:score_2<=s43[22];
							758:score_2<=s43[21];
							759:score_2<=s43[20];
							760:score_2<=s43[19];
							761:score_2<=s43[18];
							762:score_2<=s43[17];
							763:score_2<=s43[16];
							764:score_2<=s43[15];
							765:score_2<=s43[14];
							766:score_2<=s43[13];
							767:score_2<=s43[12];
							768:score_2<=s43[11];
							769:score_2<=s43[10];
							770:score_2<=s43[9];
							771:score_2<=s43[8];
							772:score_2<=s43[7];
							773:score_2<=s43[6];
							774:score_2<=s43[5];
							775:score_2<=s43[4];
							776:score_2<=s43[3];
							777:score_2<=s43[2];
							778:score_2<=s43[1];
							779:score_2<=s43[0];
							default:score_2<=0;
						endcase
					end
					592: begin
						case(col)
							730:score_2<=s42[49];
							731:score_2<=s42[48];
							732:score_2<=s42[47];
							733:score_2<=s42[46];
							734:score_2<=s42[45];
							735:score_2<=s42[44];
							736:score_2<=s42[43];
							737:score_2<=s42[42];
							738:score_2<=s42[41];
							739:score_2<=s42[40];
							740:score_2<=s42[39];
							741:score_2<=s42[38];
							742:score_2<=s42[37];
							743:score_2<=s42[36];
							744:score_2<=s42[35];
							745:score_2<=s42[34];
							746:score_2<=s42[33];
							747:score_2<=s42[32];
							748:score_2<=s42[31];
							749:score_2<=s42[30];
							750:score_2<=s42[29];
							751:score_2<=s42[28];
							752:score_2<=s42[27];
							753:score_2<=s42[26];
							754:score_2<=s42[25];
							755:score_2<=s42[24];
							756:score_2<=s42[23];
							757:score_2<=s42[22];
							758:score_2<=s42[21];
							759:score_2<=s42[20];
							760:score_2<=s42[19];
							761:score_2<=s42[18];
							762:score_2<=s42[17];
							763:score_2<=s42[16];
							764:score_2<=s42[15];
							765:score_2<=s42[14];
							766:score_2<=s42[13];
							767:score_2<=s42[12];
							768:score_2<=s42[11];
							769:score_2<=s42[10];
							770:score_2<=s42[9];
							771:score_2<=s42[8];
							772:score_2<=s42[7];
							773:score_2<=s42[6];
							774:score_2<=s42[5];
							775:score_2<=s42[4];
							776:score_2<=s42[3];
							777:score_2<=s42[2];
							778:score_2<=s42[1];
							779:score_2<=s42[0];
							default:score_2<=0;
						endcase
					end
					591: begin
						case(col)
							730:score_2<=s41[49];
							731:score_2<=s41[48];
							732:score_2<=s41[47];
							733:score_2<=s41[46];
							734:score_2<=s41[45];
							735:score_2<=s41[44];
							736:score_2<=s41[43];
							737:score_2<=s41[42];
							738:score_2<=s41[41];
							739:score_2<=s41[40];
							740:score_2<=s41[39];
							741:score_2<=s41[38];
							742:score_2<=s41[37];
							743:score_2<=s41[36];
							744:score_2<=s41[35];
							745:score_2<=s41[34];
							746:score_2<=s41[33];
							747:score_2<=s41[32];
							748:score_2<=s41[31];
							749:score_2<=s41[30];
							750:score_2<=s41[29];
							751:score_2<=s41[28];
							752:score_2<=s41[27];
							753:score_2<=s41[26];
							754:score_2<=s41[25];
							755:score_2<=s41[24];
							756:score_2<=s41[23];
							757:score_2<=s41[22];
							758:score_2<=s41[21];
							759:score_2<=s41[20];
							760:score_2<=s41[19];
							761:score_2<=s41[18];
							762:score_2<=s41[17];
							763:score_2<=s41[16];
							764:score_2<=s41[15];
							765:score_2<=s41[14];
							766:score_2<=s41[13];
							767:score_2<=s41[12];
							768:score_2<=s41[11];
							769:score_2<=s41[10];
							770:score_2<=s41[9];
							771:score_2<=s41[8];
							772:score_2<=s41[7];
							773:score_2<=s41[6];
							774:score_2<=s41[5];
							775:score_2<=s41[4];
							776:score_2<=s41[3];
							777:score_2<=s41[2];
							778:score_2<=s41[1];
							779:score_2<=s41[0];
							default:score_2<=0;
						endcase
					end
					590: begin
						case(col)
							730:score_2<=s40[49];
							731:score_2<=s40[48];
							732:score_2<=s40[47];
							733:score_2<=s40[46];
							734:score_2<=s40[45];
							735:score_2<=s40[44];
							736:score_2<=s40[43];
							737:score_2<=s40[42];
							738:score_2<=s40[41];
							739:score_2<=s40[40];
							740:score_2<=s40[39];
							741:score_2<=s40[38];
							742:score_2<=s40[37];
							743:score_2<=s40[36];
							744:score_2<=s40[35];
							745:score_2<=s40[34];
							746:score_2<=s40[33];
							747:score_2<=s40[32];
							748:score_2<=s40[31];
							749:score_2<=s40[30];
							750:score_2<=s40[29];
							751:score_2<=s40[28];
							752:score_2<=s40[27];
							753:score_2<=s40[26];
							754:score_2<=s40[25];
							755:score_2<=s40[24];
							756:score_2<=s40[23];
							757:score_2<=s40[22];
							758:score_2<=s40[21];
							759:score_2<=s40[20];
							760:score_2<=s40[19];
							761:score_2<=s40[18];
							762:score_2<=s40[17];
							763:score_2<=s40[16];
							764:score_2<=s40[15];
							765:score_2<=s40[14];
							766:score_2<=s40[13];
							767:score_2<=s40[12];
							768:score_2<=s40[11];
							769:score_2<=s40[10];
							770:score_2<=s40[9];
							771:score_2<=s40[8];
							772:score_2<=s40[7];
							773:score_2<=s40[6];
							774:score_2<=s40[5];
							775:score_2<=s40[4];
							776:score_2<=s40[3];
							777:score_2<=s40[2];
							778:score_2<=s40[1];
							779:score_2<=s40[0];
							default:score_2<=0;
						endcase
					end
					589: begin
						case(col)
							730:score_2<=s39[49];
							731:score_2<=s39[48];
							732:score_2<=s39[47];
							733:score_2<=s39[46];
							734:score_2<=s39[45];
							735:score_2<=s39[44];
							736:score_2<=s39[43];
							737:score_2<=s39[42];
							738:score_2<=s39[41];
							739:score_2<=s39[40];
							740:score_2<=s39[39];
							741:score_2<=s39[38];
							742:score_2<=s39[37];
							743:score_2<=s39[36];
							744:score_2<=s39[35];
							745:score_2<=s39[34];
							746:score_2<=s39[33];
							747:score_2<=s39[32];
							748:score_2<=s39[31];
							749:score_2<=s39[30];
							750:score_2<=s39[29];
							751:score_2<=s39[28];
							752:score_2<=s39[27];
							753:score_2<=s39[26];
							754:score_2<=s39[25];
							755:score_2<=s39[24];
							756:score_2<=s39[23];
							757:score_2<=s39[22];
							758:score_2<=s39[21];
							759:score_2<=s39[20];
							760:score_2<=s39[19];
							761:score_2<=s39[18];
							762:score_2<=s39[17];
							763:score_2<=s39[16];
							764:score_2<=s39[15];
							765:score_2<=s39[14];
							766:score_2<=s39[13];
							767:score_2<=s39[12];
							768:score_2<=s39[11];
							769:score_2<=s39[10];
							770:score_2<=s39[9];
							771:score_2<=s39[8];
							772:score_2<=s39[7];
							773:score_2<=s39[6];
							774:score_2<=s39[5];
							775:score_2<=s39[4];
							776:score_2<=s39[3];
							777:score_2<=s39[2];
							778:score_2<=s39[1];
							779:score_2<=s39[0];
							default:score_2<=0;
						endcase
					end
					588: begin
						case(col)
							730:score_2<=s38[49];
							731:score_2<=s38[48];
							732:score_2<=s38[47];
							733:score_2<=s38[46];
							734:score_2<=s38[45];
							735:score_2<=s38[44];
							736:score_2<=s38[43];
							737:score_2<=s38[42];
							738:score_2<=s38[41];
							739:score_2<=s38[40];
							740:score_2<=s38[39];
							741:score_2<=s38[38];
							742:score_2<=s38[37];
							743:score_2<=s38[36];
							744:score_2<=s38[35];
							745:score_2<=s38[34];
							746:score_2<=s38[33];
							747:score_2<=s38[32];
							748:score_2<=s38[31];
							749:score_2<=s38[30];
							750:score_2<=s38[29];
							751:score_2<=s38[28];
							752:score_2<=s38[27];
							753:score_2<=s38[26];
							754:score_2<=s38[25];
							755:score_2<=s38[24];
							756:score_2<=s38[23];
							757:score_2<=s38[22];
							758:score_2<=s38[21];
							759:score_2<=s38[20];
							760:score_2<=s38[19];
							761:score_2<=s38[18];
							762:score_2<=s38[17];
							763:score_2<=s38[16];
							764:score_2<=s38[15];
							765:score_2<=s38[14];
							766:score_2<=s38[13];
							767:score_2<=s38[12];
							768:score_2<=s38[11];
							769:score_2<=s38[10];
							770:score_2<=s38[9];
							771:score_2<=s38[8];
							772:score_2<=s38[7];
							773:score_2<=s38[6];
							774:score_2<=s38[5];
							775:score_2<=s38[4];
							776:score_2<=s38[3];
							777:score_2<=s38[2];
							778:score_2<=s38[1];
							779:score_2<=s38[0];
							default:score_2<=0;
						endcase
					end
					587: begin
						case(col)
							730:score_2<=s37[49];
							731:score_2<=s37[48];
							732:score_2<=s37[47];
							733:score_2<=s37[46];
							734:score_2<=s37[45];
							735:score_2<=s37[44];
							736:score_2<=s37[43];
							737:score_2<=s37[42];
							738:score_2<=s37[41];
							739:score_2<=s37[40];
							740:score_2<=s37[39];
							741:score_2<=s37[38];
							742:score_2<=s37[37];
							743:score_2<=s37[36];
							744:score_2<=s37[35];
							745:score_2<=s37[34];
							746:score_2<=s37[33];
							747:score_2<=s37[32];
							748:score_2<=s37[31];
							749:score_2<=s37[30];
							750:score_2<=s37[29];
							751:score_2<=s37[28];
							752:score_2<=s37[27];
							753:score_2<=s37[26];
							754:score_2<=s37[25];
							755:score_2<=s37[24];
							756:score_2<=s37[23];
							757:score_2<=s37[22];
							758:score_2<=s37[21];
							759:score_2<=s37[20];
							760:score_2<=s37[19];
							761:score_2<=s37[18];
							762:score_2<=s37[17];
							763:score_2<=s37[16];
							764:score_2<=s37[15];
							765:score_2<=s37[14];
							766:score_2<=s37[13];
							767:score_2<=s37[12];
							768:score_2<=s37[11];
							769:score_2<=s37[10];
							770:score_2<=s37[9];
							771:score_2<=s37[8];
							772:score_2<=s37[7];
							773:score_2<=s37[6];
							774:score_2<=s37[5];
							775:score_2<=s37[4];
							776:score_2<=s37[3];
							777:score_2<=s37[2];
							778:score_2<=s37[1];
							779:score_2<=s37[0];
							default:score_2<=0;
						endcase
					end
					586: begin
						case(col)
							730:score_2<=s36[49];
							731:score_2<=s36[48];
							732:score_2<=s36[47];
							733:score_2<=s36[46];
							734:score_2<=s36[45];
							735:score_2<=s36[44];
							736:score_2<=s36[43];
							737:score_2<=s36[42];
							738:score_2<=s36[41];
							739:score_2<=s36[40];
							740:score_2<=s36[39];
							741:score_2<=s36[38];
							742:score_2<=s36[37];
							743:score_2<=s36[36];
							744:score_2<=s36[35];
							745:score_2<=s36[34];
							746:score_2<=s36[33];
							747:score_2<=s36[32];
							748:score_2<=s36[31];
							749:score_2<=s36[30];
							750:score_2<=s36[29];
							751:score_2<=s36[28];
							752:score_2<=s36[27];
							753:score_2<=s36[26];
							754:score_2<=s36[25];
							755:score_2<=s36[24];
							756:score_2<=s36[23];
							757:score_2<=s36[22];
							758:score_2<=s36[21];
							759:score_2<=s36[20];
							760:score_2<=s36[19];
							761:score_2<=s36[18];
							762:score_2<=s36[17];
							763:score_2<=s36[16];
							764:score_2<=s36[15];
							765:score_2<=s36[14];
							766:score_2<=s36[13];
							767:score_2<=s36[12];
							768:score_2<=s36[11];
							769:score_2<=s36[10];
							770:score_2<=s36[9];
							771:score_2<=s36[8];
							772:score_2<=s36[7];
							773:score_2<=s36[6];
							774:score_2<=s36[5];
							775:score_2<=s36[4];
							776:score_2<=s36[3];
							777:score_2<=s36[2];
							778:score_2<=s36[1];
							779:score_2<=s36[0];
							default:score_2<=0;
						endcase
					end
					585: begin
						case(col)
							730:score_2<=s35[49];
							731:score_2<=s35[48];
							732:score_2<=s35[47];
							733:score_2<=s35[46];
							734:score_2<=s35[45];
							735:score_2<=s35[44];
							736:score_2<=s35[43];
							737:score_2<=s35[42];
							738:score_2<=s35[41];
							739:score_2<=s35[40];
							740:score_2<=s35[39];
							741:score_2<=s35[38];
							742:score_2<=s35[37];
							743:score_2<=s35[36];
							744:score_2<=s35[35];
							745:score_2<=s35[34];
							746:score_2<=s35[33];
							747:score_2<=s35[32];
							748:score_2<=s35[31];
							749:score_2<=s35[30];
							750:score_2<=s35[29];
							751:score_2<=s35[28];
							752:score_2<=s35[27];
							753:score_2<=s35[26];
							754:score_2<=s35[25];
							755:score_2<=s35[24];
							756:score_2<=s35[23];
							757:score_2<=s35[22];
							758:score_2<=s35[21];
							759:score_2<=s35[20];
							760:score_2<=s35[19];
							761:score_2<=s35[18];
							762:score_2<=s35[17];
							763:score_2<=s35[16];
							764:score_2<=s35[15];
							765:score_2<=s35[14];
							766:score_2<=s35[13];
							767:score_2<=s35[12];
							768:score_2<=s35[11];
							769:score_2<=s35[10];
							770:score_2<=s35[9];
							771:score_2<=s35[8];
							772:score_2<=s35[7];
							773:score_2<=s35[6];
							774:score_2<=s35[5];
							775:score_2<=s35[4];
							776:score_2<=s35[3];
							777:score_2<=s35[2];
							778:score_2<=s35[1];
							779:score_2<=s35[0];
							default:score_2<=0;
						endcase
					end
					584: begin
						case(col)
							730:score_2<=s34[49];
							731:score_2<=s34[48];
							732:score_2<=s34[47];
							733:score_2<=s34[46];
							734:score_2<=s34[45];
							735:score_2<=s34[44];
							736:score_2<=s34[43];
							737:score_2<=s34[42];
							738:score_2<=s34[41];
							739:score_2<=s34[40];
							740:score_2<=s34[39];
							741:score_2<=s34[38];
							742:score_2<=s34[37];
							743:score_2<=s34[36];
							744:score_2<=s34[35];
							745:score_2<=s34[34];
							746:score_2<=s34[33];
							747:score_2<=s34[32];
							748:score_2<=s34[31];
							749:score_2<=s34[30];
							750:score_2<=s34[29];
							751:score_2<=s34[28];
							752:score_2<=s34[27];
							753:score_2<=s34[26];
							754:score_2<=s34[25];
							755:score_2<=s34[24];
							756:score_2<=s34[23];
							757:score_2<=s34[22];
							758:score_2<=s34[21];
							759:score_2<=s34[20];
							760:score_2<=s34[19];
							761:score_2<=s34[18];
							762:score_2<=s34[17];
							763:score_2<=s34[16];
							764:score_2<=s34[15];
							765:score_2<=s34[14];
							766:score_2<=s34[13];
							767:score_2<=s34[12];
							768:score_2<=s34[11];
							769:score_2<=s34[10];
							770:score_2<=s34[9];
							771:score_2<=s34[8];
							772:score_2<=s34[7];
							773:score_2<=s34[6];
							774:score_2<=s34[5];
							775:score_2<=s34[4];
							776:score_2<=s34[3];
							777:score_2<=s34[2];
							778:score_2<=s34[1];
							779:score_2<=s34[0];
							default:score_2<=0;
						endcase
					end
					583: begin
						case(col)
							730:score_2<=s33[49];
							731:score_2<=s33[48];
							732:score_2<=s33[47];
							733:score_2<=s33[46];
							734:score_2<=s33[45];
							735:score_2<=s33[44];
							736:score_2<=s33[43];
							737:score_2<=s33[42];
							738:score_2<=s33[41];
							739:score_2<=s33[40];
							740:score_2<=s33[39];
							741:score_2<=s33[38];
							742:score_2<=s33[37];
							743:score_2<=s33[36];
							744:score_2<=s33[35];
							745:score_2<=s33[34];
							746:score_2<=s33[33];
							747:score_2<=s33[32];
							748:score_2<=s33[31];
							749:score_2<=s33[30];
							750:score_2<=s33[29];
							751:score_2<=s33[28];
							752:score_2<=s33[27];
							753:score_2<=s33[26];
							754:score_2<=s33[25];
							755:score_2<=s33[24];
							756:score_2<=s33[23];
							757:score_2<=s33[22];
							758:score_2<=s33[21];
							759:score_2<=s33[20];
							760:score_2<=s33[19];
							761:score_2<=s33[18];
							762:score_2<=s33[17];
							763:score_2<=s33[16];
							764:score_2<=s33[15];
							765:score_2<=s33[14];
							766:score_2<=s33[13];
							767:score_2<=s33[12];
							768:score_2<=s33[11];
							769:score_2<=s33[10];
							770:score_2<=s33[9];
							771:score_2<=s33[8];
							772:score_2<=s33[7];
							773:score_2<=s33[6];
							774:score_2<=s33[5];
							775:score_2<=s33[4];
							776:score_2<=s33[3];
							777:score_2<=s33[2];
							778:score_2<=s33[1];
							779:score_2<=s33[0];
							default:score_2<=0;
						endcase
					end
					582: begin
						case(col)
							730:score_2<=s32[49];
							731:score_2<=s32[48];
							732:score_2<=s32[47];
							733:score_2<=s32[46];
							734:score_2<=s32[45];
							735:score_2<=s32[44];
							736:score_2<=s32[43];
							737:score_2<=s32[42];
							738:score_2<=s32[41];
							739:score_2<=s32[40];
							740:score_2<=s32[39];
							741:score_2<=s32[38];
							742:score_2<=s32[37];
							743:score_2<=s32[36];
							744:score_2<=s32[35];
							745:score_2<=s32[34];
							746:score_2<=s32[33];
							747:score_2<=s32[32];
							748:score_2<=s32[31];
							749:score_2<=s32[30];
							750:score_2<=s32[29];
							751:score_2<=s32[28];
							752:score_2<=s32[27];
							753:score_2<=s32[26];
							754:score_2<=s32[25];
							755:score_2<=s32[24];
							756:score_2<=s32[23];
							757:score_2<=s32[22];
							758:score_2<=s32[21];
							759:score_2<=s32[20];
							760:score_2<=s32[19];
							761:score_2<=s32[18];
							762:score_2<=s32[17];
							763:score_2<=s32[16];
							764:score_2<=s32[15];
							765:score_2<=s32[14];
							766:score_2<=s32[13];
							767:score_2<=s32[12];
							768:score_2<=s32[11];
							769:score_2<=s32[10];
							770:score_2<=s32[9];
							771:score_2<=s32[8];
							772:score_2<=s32[7];
							773:score_2<=s32[6];
							774:score_2<=s32[5];
							775:score_2<=s32[4];
							776:score_2<=s32[3];
							777:score_2<=s32[2];
							778:score_2<=s32[1];
							779:score_2<=s32[0];
							default:score_2<=0;
						endcase
					end
					581: begin
						case(col)
							730:score_2<=s31[49];
							731:score_2<=s31[48];
							732:score_2<=s31[47];
							733:score_2<=s31[46];
							734:score_2<=s31[45];
							735:score_2<=s31[44];
							736:score_2<=s31[43];
							737:score_2<=s31[42];
							738:score_2<=s31[41];
							739:score_2<=s31[40];
							740:score_2<=s31[39];
							741:score_2<=s31[38];
							742:score_2<=s31[37];
							743:score_2<=s31[36];
							744:score_2<=s31[35];
							745:score_2<=s31[34];
							746:score_2<=s31[33];
							747:score_2<=s31[32];
							748:score_2<=s31[31];
							749:score_2<=s31[30];
							750:score_2<=s31[29];
							751:score_2<=s31[28];
							752:score_2<=s31[27];
							753:score_2<=s31[26];
							754:score_2<=s31[25];
							755:score_2<=s31[24];
							756:score_2<=s31[23];
							757:score_2<=s31[22];
							758:score_2<=s31[21];
							759:score_2<=s31[20];
							760:score_2<=s31[19];
							761:score_2<=s31[18];
							762:score_2<=s31[17];
							763:score_2<=s31[16];
							764:score_2<=s31[15];
							765:score_2<=s31[14];
							766:score_2<=s31[13];
							767:score_2<=s31[12];
							768:score_2<=s31[11];
							769:score_2<=s31[10];
							770:score_2<=s31[9];
							771:score_2<=s31[8];
							772:score_2<=s31[7];
							773:score_2<=s31[6];
							774:score_2<=s31[5];
							775:score_2<=s31[4];
							776:score_2<=s31[3];
							777:score_2<=s31[2];
							778:score_2<=s31[1];
							779:score_2<=s31[0];
							default:score_2<=0;
						endcase
					end
					580: begin
						case(col)
							730:score_2<=s30[49];
							731:score_2<=s30[48];
							732:score_2<=s30[47];
							733:score_2<=s30[46];
							734:score_2<=s30[45];
							735:score_2<=s30[44];
							736:score_2<=s30[43];
							737:score_2<=s30[42];
							738:score_2<=s30[41];
							739:score_2<=s30[40];
							740:score_2<=s30[39];
							741:score_2<=s30[38];
							742:score_2<=s30[37];
							743:score_2<=s30[36];
							744:score_2<=s30[35];
							745:score_2<=s30[34];
							746:score_2<=s30[33];
							747:score_2<=s30[32];
							748:score_2<=s30[31];
							749:score_2<=s30[30];
							750:score_2<=s30[29];
							751:score_2<=s30[28];
							752:score_2<=s30[27];
							753:score_2<=s30[26];
							754:score_2<=s30[25];
							755:score_2<=s30[24];
							756:score_2<=s30[23];
							757:score_2<=s30[22];
							758:score_2<=s30[21];
							759:score_2<=s30[20];
							760:score_2<=s30[19];
							761:score_2<=s30[18];
							762:score_2<=s30[17];
							763:score_2<=s30[16];
							764:score_2<=s30[15];
							765:score_2<=s30[14];
							766:score_2<=s30[13];
							767:score_2<=s30[12];
							768:score_2<=s30[11];
							769:score_2<=s30[10];
							770:score_2<=s30[9];
							771:score_2<=s30[8];
							772:score_2<=s30[7];
							773:score_2<=s30[6];
							774:score_2<=s30[5];
							775:score_2<=s30[4];
							776:score_2<=s30[3];
							777:score_2<=s30[2];
							778:score_2<=s30[1];
							779:score_2<=s30[0];
							default:score_2<=0;
						endcase
					end
					579: begin
						case(col)
							730:score_2<=s29[49];
							731:score_2<=s29[48];
							732:score_2<=s29[47];
							733:score_2<=s29[46];
							734:score_2<=s29[45];
							735:score_2<=s29[44];
							736:score_2<=s29[43];
							737:score_2<=s29[42];
							738:score_2<=s29[41];
							739:score_2<=s29[40];
							740:score_2<=s29[39];
							741:score_2<=s29[38];
							742:score_2<=s29[37];
							743:score_2<=s29[36];
							744:score_2<=s29[35];
							745:score_2<=s29[34];
							746:score_2<=s29[33];
							747:score_2<=s29[32];
							748:score_2<=s29[31];
							749:score_2<=s29[30];
							750:score_2<=s29[29];
							751:score_2<=s29[28];
							752:score_2<=s29[27];
							753:score_2<=s29[26];
							754:score_2<=s29[25];
							755:score_2<=s29[24];
							756:score_2<=s29[23];
							757:score_2<=s29[22];
							758:score_2<=s29[21];
							759:score_2<=s29[20];
							760:score_2<=s29[19];
							761:score_2<=s29[18];
							762:score_2<=s29[17];
							763:score_2<=s29[16];
							764:score_2<=s29[15];
							765:score_2<=s29[14];
							766:score_2<=s29[13];
							767:score_2<=s29[12];
							768:score_2<=s29[11];
							769:score_2<=s29[10];
							770:score_2<=s29[9];
							771:score_2<=s29[8];
							772:score_2<=s29[7];
							773:score_2<=s29[6];
							774:score_2<=s29[5];
							775:score_2<=s29[4];
							776:score_2<=s29[3];
							777:score_2<=s29[2];
							778:score_2<=s29[1];
							779:score_2<=s29[0];
							default:score_2<=0;
						endcase
					end
					578: begin
						case(col)
							730:score_2<=s28[49];
							731:score_2<=s28[48];
							732:score_2<=s28[47];
							733:score_2<=s28[46];
							734:score_2<=s28[45];
							735:score_2<=s28[44];
							736:score_2<=s28[43];
							737:score_2<=s28[42];
							738:score_2<=s28[41];
							739:score_2<=s28[40];
							740:score_2<=s28[39];
							741:score_2<=s28[38];
							742:score_2<=s28[37];
							743:score_2<=s28[36];
							744:score_2<=s28[35];
							745:score_2<=s28[34];
							746:score_2<=s28[33];
							747:score_2<=s28[32];
							748:score_2<=s28[31];
							749:score_2<=s28[30];
							750:score_2<=s28[29];
							751:score_2<=s28[28];
							752:score_2<=s28[27];
							753:score_2<=s28[26];
							754:score_2<=s28[25];
							755:score_2<=s28[24];
							756:score_2<=s28[23];
							757:score_2<=s28[22];
							758:score_2<=s28[21];
							759:score_2<=s28[20];
							760:score_2<=s28[19];
							761:score_2<=s28[18];
							762:score_2<=s28[17];
							763:score_2<=s28[16];
							764:score_2<=s28[15];
							765:score_2<=s28[14];
							766:score_2<=s28[13];
							767:score_2<=s28[12];
							768:score_2<=s28[11];
							769:score_2<=s28[10];
							770:score_2<=s28[9];
							771:score_2<=s28[8];
							772:score_2<=s28[7];
							773:score_2<=s28[6];
							774:score_2<=s28[5];
							775:score_2<=s28[4];
							776:score_2<=s28[3];
							777:score_2<=s28[2];
							778:score_2<=s28[1];
							779:score_2<=s28[0];
							default:score_2<=0;
						endcase
					end
					577: begin
						case(col)
							730:score_2<=s27[49];
							731:score_2<=s27[48];
							732:score_2<=s27[47];
							733:score_2<=s27[46];
							734:score_2<=s27[45];
							735:score_2<=s27[44];
							736:score_2<=s27[43];
							737:score_2<=s27[42];
							738:score_2<=s27[41];
							739:score_2<=s27[40];
							740:score_2<=s27[39];
							741:score_2<=s27[38];
							742:score_2<=s27[37];
							743:score_2<=s27[36];
							744:score_2<=s27[35];
							745:score_2<=s27[34];
							746:score_2<=s27[33];
							747:score_2<=s27[32];
							748:score_2<=s27[31];
							749:score_2<=s27[30];
							750:score_2<=s27[29];
							751:score_2<=s27[28];
							752:score_2<=s27[27];
							753:score_2<=s27[26];
							754:score_2<=s27[25];
							755:score_2<=s27[24];
							756:score_2<=s27[23];
							757:score_2<=s27[22];
							758:score_2<=s27[21];
							759:score_2<=s27[20];
							760:score_2<=s27[19];
							761:score_2<=s27[18];
							762:score_2<=s27[17];
							763:score_2<=s27[16];
							764:score_2<=s27[15];
							765:score_2<=s27[14];
							766:score_2<=s27[13];
							767:score_2<=s27[12];
							768:score_2<=s27[11];
							769:score_2<=s27[10];
							770:score_2<=s27[9];
							771:score_2<=s27[8];
							772:score_2<=s27[7];
							773:score_2<=s27[6];
							774:score_2<=s27[5];
							775:score_2<=s27[4];
							776:score_2<=s27[3];
							777:score_2<=s27[2];
							778:score_2<=s27[1];
							779:score_2<=s27[0];
							default:score_2<=0;
						endcase
					end
					576: begin
						case(col)
							730:score_2<=s26[49];
							731:score_2<=s26[48];
							732:score_2<=s26[47];
							733:score_2<=s26[46];
							734:score_2<=s26[45];
							735:score_2<=s26[44];
							736:score_2<=s26[43];
							737:score_2<=s26[42];
							738:score_2<=s26[41];
							739:score_2<=s26[40];
							740:score_2<=s26[39];
							741:score_2<=s26[38];
							742:score_2<=s26[37];
							743:score_2<=s26[36];
							744:score_2<=s26[35];
							745:score_2<=s26[34];
							746:score_2<=s26[33];
							747:score_2<=s26[32];
							748:score_2<=s26[31];
							749:score_2<=s26[30];
							750:score_2<=s26[29];
							751:score_2<=s26[28];
							752:score_2<=s26[27];
							753:score_2<=s26[26];
							754:score_2<=s26[25];
							755:score_2<=s26[24];
							756:score_2<=s26[23];
							757:score_2<=s26[22];
							758:score_2<=s26[21];
							759:score_2<=s26[20];
							760:score_2<=s26[19];
							761:score_2<=s26[18];
							762:score_2<=s26[17];
							763:score_2<=s26[16];
							764:score_2<=s26[15];
							765:score_2<=s26[14];
							766:score_2<=s26[13];
							767:score_2<=s26[12];
							768:score_2<=s26[11];
							769:score_2<=s26[10];
							770:score_2<=s26[9];
							771:score_2<=s26[8];
							772:score_2<=s26[7];
							773:score_2<=s26[6];
							774:score_2<=s26[5];
							775:score_2<=s26[4];
							776:score_2<=s26[3];
							777:score_2<=s26[2];
							778:score_2<=s26[1];
							779:score_2<=s26[0];
							default:score_2<=0;
						endcase
					end
					575: begin
						case(col)
							730:score_2<=s25[49];
							731:score_2<=s25[48];
							732:score_2<=s25[47];
							733:score_2<=s25[46];
							734:score_2<=s25[45];
							735:score_2<=s25[44];
							736:score_2<=s25[43];
							737:score_2<=s25[42];
							738:score_2<=s25[41];
							739:score_2<=s25[40];
							740:score_2<=s25[39];
							741:score_2<=s25[38];
							742:score_2<=s25[37];
							743:score_2<=s25[36];
							744:score_2<=s25[35];
							745:score_2<=s25[34];
							746:score_2<=s25[33];
							747:score_2<=s25[32];
							748:score_2<=s25[31];
							749:score_2<=s25[30];
							750:score_2<=s25[29];
							751:score_2<=s25[28];
							752:score_2<=s25[27];
							753:score_2<=s25[26];
							754:score_2<=s25[25];
							755:score_2<=s25[24];
							756:score_2<=s25[23];
							757:score_2<=s25[22];
							758:score_2<=s25[21];
							759:score_2<=s25[20];
							760:score_2<=s25[19];
							761:score_2<=s25[18];
							762:score_2<=s25[17];
							763:score_2<=s25[16];
							764:score_2<=s25[15];
							765:score_2<=s25[14];
							766:score_2<=s25[13];
							767:score_2<=s25[12];
							768:score_2<=s25[11];
							769:score_2<=s25[10];
							770:score_2<=s25[9];
							771:score_2<=s25[8];
							772:score_2<=s25[7];
							773:score_2<=s25[6];
							774:score_2<=s25[5];
							775:score_2<=s25[4];
							776:score_2<=s25[3];
							777:score_2<=s25[2];
							778:score_2<=s25[1];
							779:score_2<=s25[0];
							default:score_2<=0;
						endcase
					end
					574: begin
						case(col)
							730:score_2<=s24[49];
							731:score_2<=s24[48];
							732:score_2<=s24[47];
							733:score_2<=s24[46];
							734:score_2<=s24[45];
							735:score_2<=s24[44];
							736:score_2<=s24[43];
							737:score_2<=s24[42];
							738:score_2<=s24[41];
							739:score_2<=s24[40];
							740:score_2<=s24[39];
							741:score_2<=s24[38];
							742:score_2<=s24[37];
							743:score_2<=s24[36];
							744:score_2<=s24[35];
							745:score_2<=s24[34];
							746:score_2<=s24[33];
							747:score_2<=s24[32];
							748:score_2<=s24[31];
							749:score_2<=s24[30];
							750:score_2<=s24[29];
							751:score_2<=s24[28];
							752:score_2<=s24[27];
							753:score_2<=s24[26];
							754:score_2<=s24[25];
							755:score_2<=s24[24];
							756:score_2<=s24[23];
							757:score_2<=s24[22];
							758:score_2<=s24[21];
							759:score_2<=s24[20];
							760:score_2<=s24[19];
							761:score_2<=s24[18];
							762:score_2<=s24[17];
							763:score_2<=s24[16];
							764:score_2<=s24[15];
							765:score_2<=s24[14];
							766:score_2<=s24[13];
							767:score_2<=s24[12];
							768:score_2<=s24[11];
							769:score_2<=s24[10];
							770:score_2<=s24[9];
							771:score_2<=s24[8];
							772:score_2<=s24[7];
							773:score_2<=s24[6];
							774:score_2<=s24[5];
							775:score_2<=s24[4];
							776:score_2<=s24[3];
							777:score_2<=s24[2];
							778:score_2<=s24[1];
							779:score_2<=s24[0];
							default:score_2<=0;
						endcase
					end
					573: begin
						case(col)
							730:score_2<=s23[49];
							731:score_2<=s23[48];
							732:score_2<=s23[47];
							733:score_2<=s23[46];
							734:score_2<=s23[45];
							735:score_2<=s23[44];
							736:score_2<=s23[43];
							737:score_2<=s23[42];
							738:score_2<=s23[41];
							739:score_2<=s23[40];
							740:score_2<=s23[39];
							741:score_2<=s23[38];
							742:score_2<=s23[37];
							743:score_2<=s23[36];
							744:score_2<=s23[35];
							745:score_2<=s23[34];
							746:score_2<=s23[33];
							747:score_2<=s23[32];
							748:score_2<=s23[31];
							749:score_2<=s23[30];
							750:score_2<=s23[29];
							751:score_2<=s23[28];
							752:score_2<=s23[27];
							753:score_2<=s23[26];
							754:score_2<=s23[25];
							755:score_2<=s23[24];
							756:score_2<=s23[23];
							757:score_2<=s23[22];
							758:score_2<=s23[21];
							759:score_2<=s23[20];
							760:score_2<=s23[19];
							761:score_2<=s23[18];
							762:score_2<=s23[17];
							763:score_2<=s23[16];
							764:score_2<=s23[15];
							765:score_2<=s23[14];
							766:score_2<=s23[13];
							767:score_2<=s23[12];
							768:score_2<=s23[11];
							769:score_2<=s23[10];
							770:score_2<=s23[9];
							771:score_2<=s23[8];
							772:score_2<=s23[7];
							773:score_2<=s23[6];
							774:score_2<=s23[5];
							775:score_2<=s23[4];
							776:score_2<=s23[3];
							777:score_2<=s23[2];
							778:score_2<=s23[1];
							779:score_2<=s23[0];
							default:score_2<=0;
						endcase
					end
					572: begin
						case(col)
							730:score_2<=s22[49];
							731:score_2<=s22[48];
							732:score_2<=s22[47];
							733:score_2<=s22[46];
							734:score_2<=s22[45];
							735:score_2<=s22[44];
							736:score_2<=s22[43];
							737:score_2<=s22[42];
							738:score_2<=s22[41];
							739:score_2<=s22[40];
							740:score_2<=s22[39];
							741:score_2<=s22[38];
							742:score_2<=s22[37];
							743:score_2<=s22[36];
							744:score_2<=s22[35];
							745:score_2<=s22[34];
							746:score_2<=s22[33];
							747:score_2<=s22[32];
							748:score_2<=s22[31];
							749:score_2<=s22[30];
							750:score_2<=s22[29];
							751:score_2<=s22[28];
							752:score_2<=s22[27];
							753:score_2<=s22[26];
							754:score_2<=s22[25];
							755:score_2<=s22[24];
							756:score_2<=s22[23];
							757:score_2<=s22[22];
							758:score_2<=s22[21];
							759:score_2<=s22[20];
							760:score_2<=s22[19];
							761:score_2<=s22[18];
							762:score_2<=s22[17];
							763:score_2<=s22[16];
							764:score_2<=s22[15];
							765:score_2<=s22[14];
							766:score_2<=s22[13];
							767:score_2<=s22[12];
							768:score_2<=s22[11];
							769:score_2<=s22[10];
							770:score_2<=s22[9];
							771:score_2<=s22[8];
							772:score_2<=s22[7];
							773:score_2<=s22[6];
							774:score_2<=s22[5];
							775:score_2<=s22[4];
							776:score_2<=s22[3];
							777:score_2<=s22[2];
							778:score_2<=s22[1];
							779:score_2<=s22[0];
							default:score_2<=0;
						endcase
					end
					571: begin
						case(col)
							730:score_2<=s21[49];
							731:score_2<=s21[48];
							732:score_2<=s21[47];
							733:score_2<=s21[46];
							734:score_2<=s21[45];
							735:score_2<=s21[44];
							736:score_2<=s21[43];
							737:score_2<=s21[42];
							738:score_2<=s21[41];
							739:score_2<=s21[40];
							740:score_2<=s21[39];
							741:score_2<=s21[38];
							742:score_2<=s21[37];
							743:score_2<=s21[36];
							744:score_2<=s21[35];
							745:score_2<=s21[34];
							746:score_2<=s21[33];
							747:score_2<=s21[32];
							748:score_2<=s21[31];
							749:score_2<=s21[30];
							750:score_2<=s21[29];
							751:score_2<=s21[28];
							752:score_2<=s21[27];
							753:score_2<=s21[26];
							754:score_2<=s21[25];
							755:score_2<=s21[24];
							756:score_2<=s21[23];
							757:score_2<=s21[22];
							758:score_2<=s21[21];
							759:score_2<=s21[20];
							760:score_2<=s21[19];
							761:score_2<=s21[18];
							762:score_2<=s21[17];
							763:score_2<=s21[16];
							764:score_2<=s21[15];
							765:score_2<=s21[14];
							766:score_2<=s21[13];
							767:score_2<=s21[12];
							768:score_2<=s21[11];
							769:score_2<=s21[10];
							770:score_2<=s21[9];
							771:score_2<=s21[8];
							772:score_2<=s21[7];
							773:score_2<=s21[6];
							774:score_2<=s21[5];
							775:score_2<=s21[4];
							776:score_2<=s21[3];
							777:score_2<=s21[2];
							778:score_2<=s21[1];
							779:score_2<=s21[0];
							default:score_2<=0;
						endcase
					end
					570: begin
						case(col)
							730:score_2<=s20[49];
							731:score_2<=s20[48];
							732:score_2<=s20[47];
							733:score_2<=s20[46];
							734:score_2<=s20[45];
							735:score_2<=s20[44];
							736:score_2<=s20[43];
							737:score_2<=s20[42];
							738:score_2<=s20[41];
							739:score_2<=s20[40];
							740:score_2<=s20[39];
							741:score_2<=s20[38];
							742:score_2<=s20[37];
							743:score_2<=s20[36];
							744:score_2<=s20[35];
							745:score_2<=s20[34];
							746:score_2<=s20[33];
							747:score_2<=s20[32];
							748:score_2<=s20[31];
							749:score_2<=s20[30];
							750:score_2<=s20[29];
							751:score_2<=s20[28];
							752:score_2<=s20[27];
							753:score_2<=s20[26];
							754:score_2<=s20[25];
							755:score_2<=s20[24];
							756:score_2<=s20[23];
							757:score_2<=s20[22];
							758:score_2<=s20[21];
							759:score_2<=s20[20];
							760:score_2<=s20[19];
							761:score_2<=s20[18];
							762:score_2<=s20[17];
							763:score_2<=s20[16];
							764:score_2<=s20[15];
							765:score_2<=s20[14];
							766:score_2<=s20[13];
							767:score_2<=s20[12];
							768:score_2<=s20[11];
							769:score_2<=s20[10];
							770:score_2<=s20[9];
							771:score_2<=s20[8];
							772:score_2<=s20[7];
							773:score_2<=s20[6];
							774:score_2<=s20[5];
							775:score_2<=s20[4];
							776:score_2<=s20[3];
							777:score_2<=s20[2];
							778:score_2<=s20[1];
							779:score_2<=s20[0];
							default:score_2<=0;
						endcase
					end
					569: begin
						case(col)
							730:score_2<=s19[49];
							731:score_2<=s19[48];
							732:score_2<=s19[47];
							733:score_2<=s19[46];
							734:score_2<=s19[45];
							735:score_2<=s19[44];
							736:score_2<=s19[43];
							737:score_2<=s19[42];
							738:score_2<=s19[41];
							739:score_2<=s19[40];
							740:score_2<=s19[39];
							741:score_2<=s19[38];
							742:score_2<=s19[37];
							743:score_2<=s19[36];
							744:score_2<=s19[35];
							745:score_2<=s19[34];
							746:score_2<=s19[33];
							747:score_2<=s19[32];
							748:score_2<=s19[31];
							749:score_2<=s19[30];
							750:score_2<=s19[29];
							751:score_2<=s19[28];
							752:score_2<=s19[27];
							753:score_2<=s19[26];
							754:score_2<=s19[25];
							755:score_2<=s19[24];
							756:score_2<=s19[23];
							757:score_2<=s19[22];
							758:score_2<=s19[21];
							759:score_2<=s19[20];
							760:score_2<=s19[19];
							761:score_2<=s19[18];
							762:score_2<=s19[17];
							763:score_2<=s19[16];
							764:score_2<=s19[15];
							765:score_2<=s19[14];
							766:score_2<=s19[13];
							767:score_2<=s19[12];
							768:score_2<=s19[11];
							769:score_2<=s19[10];
							770:score_2<=s19[9];
							771:score_2<=s19[8];
							772:score_2<=s19[7];
							773:score_2<=s19[6];
							774:score_2<=s19[5];
							775:score_2<=s19[4];
							776:score_2<=s19[3];
							777:score_2<=s19[2];
							778:score_2<=s19[1];
							779:score_2<=s19[0];
							default:score_2<=0;
						endcase
					end
					568: begin
						case(col)
							730:score_2<=s18[49];
							731:score_2<=s18[48];
							732:score_2<=s18[47];
							733:score_2<=s18[46];
							734:score_2<=s18[45];
							735:score_2<=s18[44];
							736:score_2<=s18[43];
							737:score_2<=s18[42];
							738:score_2<=s18[41];
							739:score_2<=s18[40];
							740:score_2<=s18[39];
							741:score_2<=s18[38];
							742:score_2<=s18[37];
							743:score_2<=s18[36];
							744:score_2<=s18[35];
							745:score_2<=s18[34];
							746:score_2<=s18[33];
							747:score_2<=s18[32];
							748:score_2<=s18[31];
							749:score_2<=s18[30];
							750:score_2<=s18[29];
							751:score_2<=s18[28];
							752:score_2<=s18[27];
							753:score_2<=s18[26];
							754:score_2<=s18[25];
							755:score_2<=s18[24];
							756:score_2<=s18[23];
							757:score_2<=s18[22];
							758:score_2<=s18[21];
							759:score_2<=s18[20];
							760:score_2<=s18[19];
							761:score_2<=s18[18];
							762:score_2<=s18[17];
							763:score_2<=s18[16];
							764:score_2<=s18[15];
							765:score_2<=s18[14];
							766:score_2<=s18[13];
							767:score_2<=s18[12];
							768:score_2<=s18[11];
							769:score_2<=s18[10];
							770:score_2<=s18[9];
							771:score_2<=s18[8];
							772:score_2<=s18[7];
							773:score_2<=s18[6];
							774:score_2<=s18[5];
							775:score_2<=s18[4];
							776:score_2<=s18[3];
							777:score_2<=s18[2];
							778:score_2<=s18[1];
							779:score_2<=s18[0];
							default:score_2<=0;
						endcase
					end
					567: begin
						case(col)
							730:score_2<=s17[49];
							731:score_2<=s17[48];
							732:score_2<=s17[47];
							733:score_2<=s17[46];
							734:score_2<=s17[45];
							735:score_2<=s17[44];
							736:score_2<=s17[43];
							737:score_2<=s17[42];
							738:score_2<=s17[41];
							739:score_2<=s17[40];
							740:score_2<=s17[39];
							741:score_2<=s17[38];
							742:score_2<=s17[37];
							743:score_2<=s17[36];
							744:score_2<=s17[35];
							745:score_2<=s17[34];
							746:score_2<=s17[33];
							747:score_2<=s17[32];
							748:score_2<=s17[31];
							749:score_2<=s17[30];
							750:score_2<=s17[29];
							751:score_2<=s17[28];
							752:score_2<=s17[27];
							753:score_2<=s17[26];
							754:score_2<=s17[25];
							755:score_2<=s17[24];
							756:score_2<=s17[23];
							757:score_2<=s17[22];
							758:score_2<=s17[21];
							759:score_2<=s17[20];
							760:score_2<=s17[19];
							761:score_2<=s17[18];
							762:score_2<=s17[17];
							763:score_2<=s17[16];
							764:score_2<=s17[15];
							765:score_2<=s17[14];
							766:score_2<=s17[13];
							767:score_2<=s17[12];
							768:score_2<=s17[11];
							769:score_2<=s17[10];
							770:score_2<=s17[9];
							771:score_2<=s17[8];
							772:score_2<=s17[7];
							773:score_2<=s17[6];
							774:score_2<=s17[5];
							775:score_2<=s17[4];
							776:score_2<=s17[3];
							777:score_2<=s17[2];
							778:score_2<=s17[1];
							779:score_2<=s17[0];
							default:score_2<=0;
						endcase
					end
					566: begin
						case(col)
							730:score_2<=s16[49];
							731:score_2<=s16[48];
							732:score_2<=s16[47];
							733:score_2<=s16[46];
							734:score_2<=s16[45];
							735:score_2<=s16[44];
							736:score_2<=s16[43];
							737:score_2<=s16[42];
							738:score_2<=s16[41];
							739:score_2<=s16[40];
							740:score_2<=s16[39];
							741:score_2<=s16[38];
							742:score_2<=s16[37];
							743:score_2<=s16[36];
							744:score_2<=s16[35];
							745:score_2<=s16[34];
							746:score_2<=s16[33];
							747:score_2<=s16[32];
							748:score_2<=s16[31];
							749:score_2<=s16[30];
							750:score_2<=s16[29];
							751:score_2<=s16[28];
							752:score_2<=s16[27];
							753:score_2<=s16[26];
							754:score_2<=s16[25];
							755:score_2<=s16[24];
							756:score_2<=s16[23];
							757:score_2<=s16[22];
							758:score_2<=s16[21];
							759:score_2<=s16[20];
							760:score_2<=s16[19];
							761:score_2<=s16[18];
							762:score_2<=s16[17];
							763:score_2<=s16[16];
							764:score_2<=s16[15];
							765:score_2<=s16[14];
							766:score_2<=s16[13];
							767:score_2<=s16[12];
							768:score_2<=s16[11];
							769:score_2<=s16[10];
							770:score_2<=s16[9];
							771:score_2<=s16[8];
							772:score_2<=s16[7];
							773:score_2<=s16[6];
							774:score_2<=s16[5];
							775:score_2<=s16[4];
							776:score_2<=s16[3];
							777:score_2<=s16[2];
							778:score_2<=s16[1];
							779:score_2<=s16[0];
							default:score_2<=0;
						endcase
					end
					565: begin
						case(col)
							730:score_2<=s15[49];
							731:score_2<=s15[48];
							732:score_2<=s15[47];
							733:score_2<=s15[46];
							734:score_2<=s15[45];
							735:score_2<=s15[44];
							736:score_2<=s15[43];
							737:score_2<=s15[42];
							738:score_2<=s15[41];
							739:score_2<=s15[40];
							740:score_2<=s15[39];
							741:score_2<=s15[38];
							742:score_2<=s15[37];
							743:score_2<=s15[36];
							744:score_2<=s15[35];
							745:score_2<=s15[34];
							746:score_2<=s15[33];
							747:score_2<=s15[32];
							748:score_2<=s15[31];
							749:score_2<=s15[30];
							750:score_2<=s15[29];
							751:score_2<=s15[28];
							752:score_2<=s15[27];
							753:score_2<=s15[26];
							754:score_2<=s15[25];
							755:score_2<=s15[24];
							756:score_2<=s15[23];
							757:score_2<=s15[22];
							758:score_2<=s15[21];
							759:score_2<=s15[20];
							760:score_2<=s15[19];
							761:score_2<=s15[18];
							762:score_2<=s15[17];
							763:score_2<=s15[16];
							764:score_2<=s15[15];
							765:score_2<=s15[14];
							766:score_2<=s15[13];
							767:score_2<=s15[12];
							768:score_2<=s15[11];
							769:score_2<=s15[10];
							770:score_2<=s15[9];
							771:score_2<=s15[8];
							772:score_2<=s15[7];
							773:score_2<=s15[6];
							774:score_2<=s15[5];
							775:score_2<=s15[4];
							776:score_2<=s15[3];
							777:score_2<=s15[2];
							778:score_2<=s15[1];
							779:score_2<=s15[0];
							default:score_2<=0;
						endcase
					end
					564: begin
						case(col)
							730:score_2<=s14[49];
							731:score_2<=s14[48];
							732:score_2<=s14[47];
							733:score_2<=s14[46];
							734:score_2<=s14[45];
							735:score_2<=s14[44];
							736:score_2<=s14[43];
							737:score_2<=s14[42];
							738:score_2<=s14[41];
							739:score_2<=s14[40];
							740:score_2<=s14[39];
							741:score_2<=s14[38];
							742:score_2<=s14[37];
							743:score_2<=s14[36];
							744:score_2<=s14[35];
							745:score_2<=s14[34];
							746:score_2<=s14[33];
							747:score_2<=s14[32];
							748:score_2<=s14[31];
							749:score_2<=s14[30];
							750:score_2<=s14[29];
							751:score_2<=s14[28];
							752:score_2<=s14[27];
							753:score_2<=s14[26];
							754:score_2<=s14[25];
							755:score_2<=s14[24];
							756:score_2<=s14[23];
							757:score_2<=s14[22];
							758:score_2<=s14[21];
							759:score_2<=s14[20];
							760:score_2<=s14[19];
							761:score_2<=s14[18];
							762:score_2<=s14[17];
							763:score_2<=s14[16];
							764:score_2<=s14[15];
							765:score_2<=s14[14];
							766:score_2<=s14[13];
							767:score_2<=s14[12];
							768:score_2<=s14[11];
							769:score_2<=s14[10];
							770:score_2<=s14[9];
							771:score_2<=s14[8];
							772:score_2<=s14[7];
							773:score_2<=s14[6];
							774:score_2<=s14[5];
							775:score_2<=s14[4];
							776:score_2<=s14[3];
							777:score_2<=s14[2];
							778:score_2<=s14[1];
							779:score_2<=s14[0];
							default:score_2<=0;
						endcase
					end
					563: begin
						case(col)
							730:score_2<=s13[49];
							731:score_2<=s13[48];
							732:score_2<=s13[47];
							733:score_2<=s13[46];
							734:score_2<=s13[45];
							735:score_2<=s13[44];
							736:score_2<=s13[43];
							737:score_2<=s13[42];
							738:score_2<=s13[41];
							739:score_2<=s13[40];
							740:score_2<=s13[39];
							741:score_2<=s13[38];
							742:score_2<=s13[37];
							743:score_2<=s13[36];
							744:score_2<=s13[35];
							745:score_2<=s13[34];
							746:score_2<=s13[33];
							747:score_2<=s13[32];
							748:score_2<=s13[31];
							749:score_2<=s13[30];
							750:score_2<=s13[29];
							751:score_2<=s13[28];
							752:score_2<=s13[27];
							753:score_2<=s13[26];
							754:score_2<=s13[25];
							755:score_2<=s13[24];
							756:score_2<=s13[23];
							757:score_2<=s13[22];
							758:score_2<=s13[21];
							759:score_2<=s13[20];
							760:score_2<=s13[19];
							761:score_2<=s13[18];
							762:score_2<=s13[17];
							763:score_2<=s13[16];
							764:score_2<=s13[15];
							765:score_2<=s13[14];
							766:score_2<=s13[13];
							767:score_2<=s13[12];
							768:score_2<=s13[11];
							769:score_2<=s13[10];
							770:score_2<=s13[9];
							771:score_2<=s13[8];
							772:score_2<=s13[7];
							773:score_2<=s13[6];
							774:score_2<=s13[5];
							775:score_2<=s13[4];
							776:score_2<=s13[3];
							777:score_2<=s13[2];
							778:score_2<=s13[1];
							779:score_2<=s13[0];
							default:score_2<=0;
						endcase
					end
					562: begin
						case(col)
							730:score_2<=s12[49];
							731:score_2<=s12[48];
							732:score_2<=s12[47];
							733:score_2<=s12[46];
							734:score_2<=s12[45];
							735:score_2<=s12[44];
							736:score_2<=s12[43];
							737:score_2<=s12[42];
							738:score_2<=s12[41];
							739:score_2<=s12[40];
							740:score_2<=s12[39];
							741:score_2<=s12[38];
							742:score_2<=s12[37];
							743:score_2<=s12[36];
							744:score_2<=s12[35];
							745:score_2<=s12[34];
							746:score_2<=s12[33];
							747:score_2<=s12[32];
							748:score_2<=s12[31];
							749:score_2<=s12[30];
							750:score_2<=s12[29];
							751:score_2<=s12[28];
							752:score_2<=s12[27];
							753:score_2<=s12[26];
							754:score_2<=s12[25];
							755:score_2<=s12[24];
							756:score_2<=s12[23];
							757:score_2<=s12[22];
							758:score_2<=s12[21];
							759:score_2<=s12[20];
							760:score_2<=s12[19];
							761:score_2<=s12[18];
							762:score_2<=s12[17];
							763:score_2<=s12[16];
							764:score_2<=s12[15];
							765:score_2<=s12[14];
							766:score_2<=s12[13];
							767:score_2<=s12[12];
							768:score_2<=s12[11];
							769:score_2<=s12[10];
							770:score_2<=s12[9];
							771:score_2<=s12[8];
							772:score_2<=s12[7];
							773:score_2<=s12[6];
							774:score_2<=s12[5];
							775:score_2<=s12[4];
							776:score_2<=s12[3];
							777:score_2<=s12[2];
							778:score_2<=s12[1];
							779:score_2<=s12[0];
							default:score_2<=0;
						endcase
					end
					561: begin
						case(col)
							730:score_2<=s11[49];
							731:score_2<=s11[48];
							732:score_2<=s11[47];
							733:score_2<=s11[46];
							734:score_2<=s11[45];
							735:score_2<=s11[44];
							736:score_2<=s11[43];
							737:score_2<=s11[42];
							738:score_2<=s11[41];
							739:score_2<=s11[40];
							740:score_2<=s11[39];
							741:score_2<=s11[38];
							742:score_2<=s11[37];
							743:score_2<=s11[36];
							744:score_2<=s11[35];
							745:score_2<=s11[34];
							746:score_2<=s11[33];
							747:score_2<=s11[32];
							748:score_2<=s11[31];
							749:score_2<=s11[30];
							750:score_2<=s11[29];
							751:score_2<=s11[28];
							752:score_2<=s11[27];
							753:score_2<=s11[26];
							754:score_2<=s11[25];
							755:score_2<=s11[24];
							756:score_2<=s11[23];
							757:score_2<=s11[22];
							758:score_2<=s11[21];
							759:score_2<=s11[20];
							760:score_2<=s11[19];
							761:score_2<=s11[18];
							762:score_2<=s11[17];
							763:score_2<=s11[16];
							764:score_2<=s11[15];
							765:score_2<=s11[14];
							766:score_2<=s11[13];
							767:score_2<=s11[12];
							768:score_2<=s11[11];
							769:score_2<=s11[10];
							770:score_2<=s11[9];
							771:score_2<=s11[8];
							772:score_2<=s11[7];
							773:score_2<=s11[6];
							774:score_2<=s11[5];
							775:score_2<=s11[4];
							776:score_2<=s11[3];
							777:score_2<=s11[2];
							778:score_2<=s11[1];
							779:score_2<=s11[0];
							default:score_2<=0;
						endcase
					end
					560: begin
						case(col)
							730:score_2<=s10[49];
							731:score_2<=s10[48];
							732:score_2<=s10[47];
							733:score_2<=s10[46];
							734:score_2<=s10[45];
							735:score_2<=s10[44];
							736:score_2<=s10[43];
							737:score_2<=s10[42];
							738:score_2<=s10[41];
							739:score_2<=s10[40];
							740:score_2<=s10[39];
							741:score_2<=s10[38];
							742:score_2<=s10[37];
							743:score_2<=s10[36];
							744:score_2<=s10[35];
							745:score_2<=s10[34];
							746:score_2<=s10[33];
							747:score_2<=s10[32];
							748:score_2<=s10[31];
							749:score_2<=s10[30];
							750:score_2<=s10[29];
							751:score_2<=s10[28];
							752:score_2<=s10[27];
							753:score_2<=s10[26];
							754:score_2<=s10[25];
							755:score_2<=s10[24];
							756:score_2<=s10[23];
							757:score_2<=s10[22];
							758:score_2<=s10[21];
							759:score_2<=s10[20];
							760:score_2<=s10[19];
							761:score_2<=s10[18];
							762:score_2<=s10[17];
							763:score_2<=s10[16];
							764:score_2<=s10[15];
							765:score_2<=s10[14];
							766:score_2<=s10[13];
							767:score_2<=s10[12];
							768:score_2<=s10[11];
							769:score_2<=s10[10];
							770:score_2<=s10[9];
							771:score_2<=s10[8];
							772:score_2<=s10[7];
							773:score_2<=s10[6];
							774:score_2<=s10[5];
							775:score_2<=s10[4];
							776:score_2<=s10[3];
							777:score_2<=s10[2];
							778:score_2<=s10[1];
							779:score_2<=s10[0];
							default:score_2<=0;
						endcase
					end
					559: begin
						case(col)
							730:score_2<=s9[49];
							731:score_2<=s9[48];
							732:score_2<=s9[47];
							733:score_2<=s9[46];
							734:score_2<=s9[45];
							735:score_2<=s9[44];
							736:score_2<=s9[43];
							737:score_2<=s9[42];
							738:score_2<=s9[41];
							739:score_2<=s9[40];
							740:score_2<=s9[39];
							741:score_2<=s9[38];
							742:score_2<=s9[37];
							743:score_2<=s9[36];
							744:score_2<=s9[35];
							745:score_2<=s9[34];
							746:score_2<=s9[33];
							747:score_2<=s9[32];
							748:score_2<=s9[31];
							749:score_2<=s9[30];
							750:score_2<=s9[29];
							751:score_2<=s9[28];
							752:score_2<=s9[27];
							753:score_2<=s9[26];
							754:score_2<=s9[25];
							755:score_2<=s9[24];
							756:score_2<=s9[23];
							757:score_2<=s9[22];
							758:score_2<=s9[21];
							759:score_2<=s9[20];
							760:score_2<=s9[19];
							761:score_2<=s9[18];
							762:score_2<=s9[17];
							763:score_2<=s9[16];
							764:score_2<=s9[15];
							765:score_2<=s9[14];
							766:score_2<=s9[13];
							767:score_2<=s9[12];
							768:score_2<=s9[11];
							769:score_2<=s9[10];
							770:score_2<=s9[9];
							771:score_2<=s9[8];
							772:score_2<=s9[7];
							773:score_2<=s9[6];
							774:score_2<=s9[5];
							775:score_2<=s9[4];
							776:score_2<=s9[3];
							777:score_2<=s9[2];
							778:score_2<=s9[1];
							779:score_2<=s9[0];
							default:score_2<=0;
						endcase
					end
					558: begin
						case(col)
							730:score_2<=s8[49];
							731:score_2<=s8[48];
							732:score_2<=s8[47];
							733:score_2<=s8[46];
							734:score_2<=s8[45];
							735:score_2<=s8[44];
							736:score_2<=s8[43];
							737:score_2<=s8[42];
							738:score_2<=s8[41];
							739:score_2<=s8[40];
							740:score_2<=s8[39];
							741:score_2<=s8[38];
							742:score_2<=s8[37];
							743:score_2<=s8[36];
							744:score_2<=s8[35];
							745:score_2<=s8[34];
							746:score_2<=s8[33];
							747:score_2<=s8[32];
							748:score_2<=s8[31];
							749:score_2<=s8[30];
							750:score_2<=s8[29];
							751:score_2<=s8[28];
							752:score_2<=s8[27];
							753:score_2<=s8[26];
							754:score_2<=s8[25];
							755:score_2<=s8[24];
							756:score_2<=s8[23];
							757:score_2<=s8[22];
							758:score_2<=s8[21];
							759:score_2<=s8[20];
							760:score_2<=s8[19];
							761:score_2<=s8[18];
							762:score_2<=s8[17];
							763:score_2<=s8[16];
							764:score_2<=s8[15];
							765:score_2<=s8[14];
							766:score_2<=s8[13];
							767:score_2<=s8[12];
							768:score_2<=s8[11];
							769:score_2<=s8[10];
							770:score_2<=s8[9];
							771:score_2<=s8[8];
							772:score_2<=s8[7];
							773:score_2<=s8[6];
							774:score_2<=s8[5];
							775:score_2<=s8[4];
							776:score_2<=s8[3];
							777:score_2<=s8[2];
							778:score_2<=s8[1];
							779:score_2<=s8[0];
							default:score_2<=0;
						endcase
					end
					557: begin
						case(col)
							730:score_2<=s7[49];
							731:score_2<=s7[48];
							732:score_2<=s7[47];
							733:score_2<=s7[46];
							734:score_2<=s7[45];
							735:score_2<=s7[44];
							736:score_2<=s7[43];
							737:score_2<=s7[42];
							738:score_2<=s7[41];
							739:score_2<=s7[40];
							740:score_2<=s7[39];
							741:score_2<=s7[38];
							742:score_2<=s7[37];
							743:score_2<=s7[36];
							744:score_2<=s7[35];
							745:score_2<=s7[34];
							746:score_2<=s7[33];
							747:score_2<=s7[32];
							748:score_2<=s7[31];
							749:score_2<=s7[30];
							750:score_2<=s7[29];
							751:score_2<=s7[28];
							752:score_2<=s7[27];
							753:score_2<=s7[26];
							754:score_2<=s7[25];
							755:score_2<=s7[24];
							756:score_2<=s7[23];
							757:score_2<=s7[22];
							758:score_2<=s7[21];
							759:score_2<=s7[20];
							760:score_2<=s7[19];
							761:score_2<=s7[18];
							762:score_2<=s7[17];
							763:score_2<=s7[16];
							764:score_2<=s7[15];
							765:score_2<=s7[14];
							766:score_2<=s7[13];
							767:score_2<=s7[12];
							768:score_2<=s7[11];
							769:score_2<=s7[10];
							770:score_2<=s7[9];
							771:score_2<=s7[8];
							772:score_2<=s7[7];
							773:score_2<=s7[6];
							774:score_2<=s7[5];
							775:score_2<=s7[4];
							776:score_2<=s7[3];
							777:score_2<=s7[2];
							778:score_2<=s7[1];
							779:score_2<=s7[0];
							default:score_2<=0;
						endcase
					end
					556: begin
						case(col)
							730:score_2<=s6[49];
							731:score_2<=s6[48];
							732:score_2<=s6[47];
							733:score_2<=s6[46];
							734:score_2<=s6[45];
							735:score_2<=s6[44];
							736:score_2<=s6[43];
							737:score_2<=s6[42];
							738:score_2<=s6[41];
							739:score_2<=s6[40];
							740:score_2<=s6[39];
							741:score_2<=s6[38];
							742:score_2<=s6[37];
							743:score_2<=s6[36];
							744:score_2<=s6[35];
							745:score_2<=s6[34];
							746:score_2<=s6[33];
							747:score_2<=s6[32];
							748:score_2<=s6[31];
							749:score_2<=s6[30];
							750:score_2<=s6[29];
							751:score_2<=s6[28];
							752:score_2<=s6[27];
							753:score_2<=s6[26];
							754:score_2<=s6[25];
							755:score_2<=s6[24];
							756:score_2<=s6[23];
							757:score_2<=s6[22];
							758:score_2<=s6[21];
							759:score_2<=s6[20];
							760:score_2<=s6[19];
							761:score_2<=s6[18];
							762:score_2<=s6[17];
							763:score_2<=s6[16];
							764:score_2<=s6[15];
							765:score_2<=s6[14];
							766:score_2<=s6[13];
							767:score_2<=s6[12];
							768:score_2<=s6[11];
							769:score_2<=s6[10];
							770:score_2<=s6[9];
							771:score_2<=s6[8];
							772:score_2<=s6[7];
							773:score_2<=s6[6];
							774:score_2<=s6[5];
							775:score_2<=s6[4];
							776:score_2<=s6[3];
							777:score_2<=s6[2];
							778:score_2<=s6[1];
							779:score_2<=s6[0];
							default:score_2<=0;
						endcase
					end
					555: begin
						case(col)
							730:score_2<=s5[49];
							731:score_2<=s5[48];
							732:score_2<=s5[47];
							733:score_2<=s5[46];
							734:score_2<=s5[45];
							735:score_2<=s5[44];
							736:score_2<=s5[43];
							737:score_2<=s5[42];
							738:score_2<=s5[41];
							739:score_2<=s5[40];
							740:score_2<=s5[39];
							741:score_2<=s5[38];
							742:score_2<=s5[37];
							743:score_2<=s5[36];
							744:score_2<=s5[35];
							745:score_2<=s5[34];
							746:score_2<=s5[33];
							747:score_2<=s5[32];
							748:score_2<=s5[31];
							749:score_2<=s5[30];
							750:score_2<=s5[29];
							751:score_2<=s5[28];
							752:score_2<=s5[27];
							753:score_2<=s5[26];
							754:score_2<=s5[25];
							755:score_2<=s5[24];
							756:score_2<=s5[23];
							757:score_2<=s5[22];
							758:score_2<=s5[21];
							759:score_2<=s5[20];
							760:score_2<=s5[19];
							761:score_2<=s5[18];
							762:score_2<=s5[17];
							763:score_2<=s5[16];
							764:score_2<=s5[15];
							765:score_2<=s5[14];
							766:score_2<=s5[13];
							767:score_2<=s5[12];
							768:score_2<=s5[11];
							769:score_2<=s5[10];
							770:score_2<=s5[9];
							771:score_2<=s5[8];
							772:score_2<=s5[7];
							773:score_2<=s5[6];
							774:score_2<=s5[5];
							775:score_2<=s5[4];
							776:score_2<=s5[3];
							777:score_2<=s5[2];
							778:score_2<=s5[1];
							779:score_2<=s5[0];
							default:score_2<=0;
						endcase
					end
					554: begin
						case(col)
							730:score_2<=s4[49];
							731:score_2<=s4[48];
							732:score_2<=s4[47];
							733:score_2<=s4[46];
							734:score_2<=s4[45];
							735:score_2<=s4[44];
							736:score_2<=s4[43];
							737:score_2<=s4[42];
							738:score_2<=s4[41];
							739:score_2<=s4[40];
							740:score_2<=s4[39];
							741:score_2<=s4[38];
							742:score_2<=s4[37];
							743:score_2<=s4[36];
							744:score_2<=s4[35];
							745:score_2<=s4[34];
							746:score_2<=s4[33];
							747:score_2<=s4[32];
							748:score_2<=s4[31];
							749:score_2<=s4[30];
							750:score_2<=s4[29];
							751:score_2<=s4[28];
							752:score_2<=s4[27];
							753:score_2<=s4[26];
							754:score_2<=s4[25];
							755:score_2<=s4[24];
							756:score_2<=s4[23];
							757:score_2<=s4[22];
							758:score_2<=s4[21];
							759:score_2<=s4[20];
							760:score_2<=s4[19];
							761:score_2<=s4[18];
							762:score_2<=s4[17];
							763:score_2<=s4[16];
							764:score_2<=s4[15];
							765:score_2<=s4[14];
							766:score_2<=s4[13];
							767:score_2<=s4[12];
							768:score_2<=s4[11];
							769:score_2<=s4[10];
							770:score_2<=s4[9];
							771:score_2<=s4[8];
							772:score_2<=s4[7];
							773:score_2<=s4[6];
							774:score_2<=s4[5];
							775:score_2<=s4[4];
							776:score_2<=s4[3];
							777:score_2<=s4[2];
							778:score_2<=s4[1];
							779:score_2<=s4[0];
							default:score_2<=0;
						endcase
					end
					553: begin
						case(col)
							730:score_2<=s3[49];
							731:score_2<=s3[48];
							732:score_2<=s3[47];
							733:score_2<=s3[46];
							734:score_2<=s3[45];
							735:score_2<=s3[44];
							736:score_2<=s3[43];
							737:score_2<=s3[42];
							738:score_2<=s3[41];
							739:score_2<=s3[40];
							740:score_2<=s3[39];
							741:score_2<=s3[38];
							742:score_2<=s3[37];
							743:score_2<=s3[36];
							744:score_2<=s3[35];
							745:score_2<=s3[34];
							746:score_2<=s3[33];
							747:score_2<=s3[32];
							748:score_2<=s3[31];
							749:score_2<=s3[30];
							750:score_2<=s3[29];
							751:score_2<=s3[28];
							752:score_2<=s3[27];
							753:score_2<=s3[26];
							754:score_2<=s3[25];
							755:score_2<=s3[24];
							756:score_2<=s3[23];
							757:score_2<=s3[22];
							758:score_2<=s3[21];
							759:score_2<=s3[20];
							760:score_2<=s3[19];
							761:score_2<=s3[18];
							762:score_2<=s3[17];
							763:score_2<=s3[16];
							764:score_2<=s3[15];
							765:score_2<=s3[14];
							766:score_2<=s3[13];
							767:score_2<=s3[12];
							768:score_2<=s3[11];
							769:score_2<=s3[10];
							770:score_2<=s3[9];
							771:score_2<=s3[8];
							772:score_2<=s3[7];
							773:score_2<=s3[6];
							774:score_2<=s3[5];
							775:score_2<=s3[4];
							776:score_2<=s3[3];
							777:score_2<=s3[2];
							778:score_2<=s3[1];
							779:score_2<=s3[0];
							default:score_2<=0;
						endcase
					end
					552: begin
						case(col)
							730:score_2<=s2[49];
							731:score_2<=s2[48];
							732:score_2<=s2[47];
							733:score_2<=s2[46];
							734:score_2<=s2[45];
							735:score_2<=s2[44];
							736:score_2<=s2[43];
							737:score_2<=s2[42];
							738:score_2<=s2[41];
							739:score_2<=s2[40];
							740:score_2<=s2[39];
							741:score_2<=s2[38];
							742:score_2<=s2[37];
							743:score_2<=s2[36];
							744:score_2<=s2[35];
							745:score_2<=s2[34];
							746:score_2<=s2[33];
							747:score_2<=s2[32];
							748:score_2<=s2[31];
							749:score_2<=s2[30];
							750:score_2<=s2[29];
							751:score_2<=s2[28];
							752:score_2<=s2[27];
							753:score_2<=s2[26];
							754:score_2<=s2[25];
							755:score_2<=s2[24];
							756:score_2<=s2[23];
							757:score_2<=s2[22];
							758:score_2<=s2[21];
							759:score_2<=s2[20];
							760:score_2<=s2[19];
							761:score_2<=s2[18];
							762:score_2<=s2[17];
							763:score_2<=s2[16];
							764:score_2<=s2[15];
							765:score_2<=s2[14];
							766:score_2<=s2[13];
							767:score_2<=s2[12];
							768:score_2<=s2[11];
							769:score_2<=s2[10];
							770:score_2<=s2[9];
							771:score_2<=s2[8];
							772:score_2<=s2[7];
							773:score_2<=s2[6];
							774:score_2<=s2[5];
							775:score_2<=s2[4];
							776:score_2<=s2[3];
							777:score_2<=s2[2];
							778:score_2<=s2[1];
							779:score_2<=s2[0];
							default:score_2<=0;
						endcase
					end
					551: begin
						case(col)
							730:score_2<=s1[49];
							731:score_2<=s1[48];
							732:score_2<=s1[47];
							733:score_2<=s1[46];
							734:score_2<=s1[45];
							735:score_2<=s1[44];
							736:score_2<=s1[43];
							737:score_2<=s1[42];
							738:score_2<=s1[41];
							739:score_2<=s1[40];
							740:score_2<=s1[39];
							741:score_2<=s1[38];
							742:score_2<=s1[37];
							743:score_2<=s1[36];
							744:score_2<=s1[35];
							745:score_2<=s1[34];
							746:score_2<=s1[33];
							747:score_2<=s1[32];
							748:score_2<=s1[31];
							749:score_2<=s1[30];
							750:score_2<=s1[29];
							751:score_2<=s1[28];
							752:score_2<=s1[27];
							753:score_2<=s1[26];
							754:score_2<=s1[25];
							755:score_2<=s1[24];
							756:score_2<=s1[23];
							757:score_2<=s1[22];
							758:score_2<=s1[21];
							759:score_2<=s1[20];
							760:score_2<=s1[19];
							761:score_2<=s1[18];
							762:score_2<=s1[17];
							763:score_2<=s1[16];
							764:score_2<=s1[15];
							765:score_2<=s1[14];
							766:score_2<=s1[13];
							767:score_2<=s1[12];
							768:score_2<=s1[11];
							769:score_2<=s1[10];
							770:score_2<=s1[9];
							771:score_2<=s1[8];
							772:score_2<=s1[7];
							773:score_2<=s1[6];
							774:score_2<=s1[5];
							775:score_2<=s1[4];
							776:score_2<=s1[3];
							777:score_2<=s1[2];
							778:score_2<=s1[1];
							779:score_2<=s1[0];
							default:score_2<=0;
						endcase
					end
			default:score_2<=0;
	endcase
end

endmodule